magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 731 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 165 47 195 177
rect 267 93 297 177
rect 455 47 485 177
rect 551 47 581 177
rect 623 47 653 177
<< scpmoshvt >>
rect 79 297 109 497
rect 165 297 195 497
rect 267 297 297 381
rect 455 297 485 497
rect 539 297 569 497
rect 623 297 653 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 165 177
rect 109 131 120 165
rect 154 131 165 165
rect 109 97 165 131
rect 109 63 120 97
rect 154 63 165 97
rect 109 47 165 63
rect 195 157 267 177
rect 195 123 206 157
rect 240 123 267 157
rect 195 93 267 123
rect 297 165 349 177
rect 297 131 307 165
rect 341 131 349 165
rect 297 93 349 131
rect 403 93 455 177
rect 195 89 252 93
rect 195 55 206 89
rect 240 55 252 89
rect 195 47 252 55
rect 403 59 411 93
rect 445 59 455 93
rect 403 47 455 59
rect 485 163 551 177
rect 485 129 498 163
rect 532 129 551 163
rect 485 47 551 129
rect 581 47 623 177
rect 653 165 705 177
rect 653 131 663 165
rect 697 131 705 165
rect 653 47 705 131
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 297 79 451
rect 109 469 165 497
rect 109 435 120 469
rect 154 435 165 469
rect 109 401 165 435
rect 109 367 120 401
rect 154 367 165 401
rect 109 297 165 367
rect 195 489 282 497
rect 195 455 224 489
rect 258 455 282 489
rect 195 435 282 455
rect 403 439 455 497
rect 195 381 252 435
rect 403 405 411 439
rect 445 405 455 439
rect 195 297 267 381
rect 297 345 349 381
rect 297 311 307 345
rect 341 311 349 345
rect 297 297 349 311
rect 403 371 455 405
rect 403 337 411 371
rect 445 337 455 371
rect 403 297 455 337
rect 485 485 539 497
rect 485 451 495 485
rect 529 451 539 485
rect 485 417 539 451
rect 485 383 495 417
rect 529 383 539 417
rect 485 297 539 383
rect 569 489 623 497
rect 569 455 579 489
rect 613 455 623 489
rect 569 297 623 455
rect 653 485 705 497
rect 653 451 663 485
rect 697 451 705 485
rect 653 417 705 451
rect 653 383 663 417
rect 697 383 705 417
rect 653 297 705 383
<< ndiffc >>
rect 35 59 69 93
rect 120 131 154 165
rect 120 63 154 97
rect 206 123 240 157
rect 307 131 341 165
rect 206 55 240 89
rect 411 59 445 93
rect 498 129 532 163
rect 663 131 697 165
<< pdiffc >>
rect 35 451 69 485
rect 120 435 154 469
rect 120 367 154 401
rect 224 455 258 489
rect 411 405 445 439
rect 307 311 341 345
rect 411 337 445 371
rect 495 451 529 485
rect 495 383 529 417
rect 579 455 613 489
rect 663 451 697 485
rect 663 383 697 417
<< poly >>
rect 79 497 109 523
rect 165 497 195 523
rect 455 497 485 523
rect 539 497 569 523
rect 623 497 653 523
rect 267 381 297 407
rect 79 259 109 297
rect 165 259 195 297
rect 267 265 297 297
rect 455 265 485 297
rect 539 265 569 297
rect 623 265 653 297
rect 79 249 195 259
rect 79 215 130 249
rect 164 215 195 249
rect 79 205 195 215
rect 79 177 109 205
rect 165 177 195 205
rect 261 249 315 265
rect 261 215 271 249
rect 305 215 315 249
rect 261 199 315 215
rect 391 249 485 265
rect 391 215 401 249
rect 435 215 485 249
rect 267 177 297 199
rect 391 198 485 215
rect 527 249 581 265
rect 527 215 537 249
rect 571 215 581 249
rect 527 199 581 215
rect 455 177 485 198
rect 551 177 581 199
rect 623 249 698 265
rect 623 215 654 249
rect 688 215 698 249
rect 623 199 698 215
rect 623 177 653 199
rect 267 67 297 93
rect 79 21 109 47
rect 165 21 195 47
rect 455 21 485 47
rect 551 21 581 47
rect 623 21 653 47
<< polycont >>
rect 130 215 164 249
rect 271 215 305 249
rect 401 215 435 249
rect 537 215 571 249
rect 654 215 688 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 485 85 527
rect 208 489 274 527
rect 18 451 35 485
rect 69 451 85 485
rect 119 469 170 485
rect 119 435 120 469
rect 154 435 170 469
rect 208 455 224 489
rect 258 455 274 489
rect 119 401 170 435
rect 395 439 445 493
rect 395 421 411 439
rect 30 367 120 401
rect 154 367 170 401
rect 223 405 411 421
rect 223 379 445 405
rect 30 177 76 367
rect 223 333 257 379
rect 411 371 445 379
rect 114 299 257 333
rect 291 311 307 345
rect 341 311 373 345
rect 114 249 180 299
rect 339 265 373 311
rect 479 485 545 493
rect 479 451 495 485
rect 529 451 545 485
rect 479 417 545 451
rect 579 489 613 527
rect 579 437 613 455
rect 647 485 713 493
rect 647 451 663 485
rect 697 451 713 485
rect 479 383 495 417
rect 529 403 545 417
rect 647 417 713 451
rect 647 403 663 417
rect 529 383 663 403
rect 697 383 713 417
rect 479 369 713 383
rect 411 335 445 337
rect 411 301 503 335
rect 114 215 130 249
rect 164 215 180 249
rect 214 249 305 265
rect 214 215 271 249
rect 214 207 305 215
rect 266 199 305 207
rect 339 249 435 265
rect 339 215 401 249
rect 339 199 435 215
rect 30 165 170 177
rect 30 143 120 165
rect 104 131 120 143
rect 154 131 170 165
rect 18 93 69 109
rect 18 59 35 93
rect 104 97 170 131
rect 104 63 120 97
rect 154 63 170 97
rect 204 157 244 173
rect 339 165 373 199
rect 204 123 206 157
rect 240 123 244 157
rect 291 131 307 165
rect 341 131 373 165
rect 469 165 503 301
rect 537 249 620 323
rect 571 215 620 249
rect 537 199 620 215
rect 654 249 712 323
rect 688 215 712 249
rect 654 199 712 215
rect 469 163 548 165
rect 469 129 498 163
rect 532 129 548 163
rect 469 127 548 129
rect 647 131 663 165
rect 697 131 713 165
rect 204 89 244 123
rect 18 17 69 59
rect 204 55 206 89
rect 240 55 244 89
rect 204 17 244 55
rect 395 59 411 93
rect 445 59 461 93
rect 395 17 461 59
rect 647 17 713 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 214 221 248 255 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 30 357 64 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 586 289 620 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a21bo_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3990100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3983804
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
