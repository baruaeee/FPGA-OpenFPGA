magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 130 582
<< pwell >>
rect 28 -11 52 11
<< obsli1 >>
rect 0 527 29 561
rect 63 527 92 561
rect 0 -17 29 17
rect 63 -17 92 17
<< obsli1c >>
rect 29 527 63 561
rect 29 -17 63 17
<< metal1 >>
rect 0 561 92 592
rect 0 527 29 561
rect 63 527 92 561
rect 0 496 92 527
rect 0 17 92 48
rect 0 -17 29 17
rect 63 -17 92 17
rect 0 -48 92 -17
<< labels >>
rlabel metal1 s 0 -48 92 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel pwell s 28 -11 52 11 8 VNB
port 2 nsew ground bidirectional
rlabel nwell s -38 261 130 582 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 496 92 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 92 544
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2152956
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2151728
<< end >>
