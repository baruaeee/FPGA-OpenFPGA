# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__corner_bus_overlay
  CLASS PAD ;
  ORIGIN  0.000000  0.000000 ;
  FOREIGN sky130_fd_io__corner_bus_overlay  0.000000  0.000000 ;
  SIZE 200 BY  203.6650 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 56.790000  0.500000 59.770000 ;
        RECT 53.125000  0.000000 56.105000  0.500000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT  0.000000 52.030000  0.575000 55.010000 ;
        RECT 48.365000  0.000000 51.345000  0.575000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.550000 1.270000 17.200000 ;
      LAYER met4 ;
        RECT 8.885000 0.000000 13.535000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 12.650000 1.270000 17.100000 ;
      LAYER met5 ;
        RECT 8.985000 0.000000 13.435000 1.270000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 5.700000 1.270000 11.150000 ;
      LAYER met4 ;
        RECT 2.035000 0.000000 7.485000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 5.800000 1.270000 11.050000 ;
      LAYER met5 ;
        RECT 2.135000 0.000000 7.385000 1.270000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 18.600000 1.255000 22.050000 ;
      LAYER met4 ;
        RECT 14.935000 0.000000 18.385000 1.255000 ;
      LAYER met5 ;
        RECT 0.000000 18.700000 1.255000 21.950000 ;
      LAYER met5 ;
        RECT 15.035000 0.000000 18.285000 1.255000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 23.450000 1.270000 28.100000 ;
      LAYER met4 ;
        RECT 0.000000 73.705000 1.270000 98.665000 ;
      LAYER met4 ;
        RECT 19.785000 0.000000 24.435000 1.270000 ;
        RECT 70.040000 0.000000 95.000000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 23.550000 1.270000 28.000000 ;
        RECT 0.000000 73.700000 1.270000 98.650000 ;
      LAYER met5 ;
        RECT 19.885000 0.000000 24.335000 1.270000 ;
        RECT 70.035000 0.000000 94.985000 1.270000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 67.750000 1.270000 72.200000 ;
      LAYER met4 ;
        RECT 64.085000 0.000000 68.535000 1.270000 ;
      LAYER met5 ;
        RECT  0.000000 67.850000  1.270000 72.100000 ;
        RECT 64.185000  0.000000 68.435000  1.270000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 40.400000 1.270000 43.850000 ;
      LAYER met4 ;
        RECT 0.000000 51.400000 1.270000 51.730000 ;
        RECT 0.000000 55.310000 1.270000 56.490000 ;
        RECT 0.000000 60.070000 1.270000 60.400000 ;
      LAYER met4 ;
        RECT 36.735000 0.000000 40.185000 1.270000 ;
        RECT 47.735000 0.000000 48.065000 1.270000 ;
        RECT 51.645000 0.000000 52.825000 1.270000 ;
        RECT 56.405000 0.000000 56.735000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 40.505000 1.270000 43.750000 ;
      LAYER met5 ;
        RECT 0.000000 51.400000 1.270000 60.400000 ;
      LAYER met5 ;
        RECT 36.840000 0.000000 40.085000 1.270000 ;
        RECT 47.735000 0.000000 56.735000 1.270000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 45.250000 1.270000 49.900000 ;
      LAYER met4 ;
        RECT 41.585000 0.000000 46.235000 1.270000 ;
      LAYER met5 ;
        RECT  0.000000 45.350000  1.270000 49.800000 ;
        RECT 41.685000  0.000000 46.135000  1.270000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT  25.835000 0.000000  30.485000 1.270000 ;
        RECT 175.785000 0.000000 200.000000 1.270000 ;
      LAYER met4 ;
        RECT 0.000000 179.450000 1.270000 203.665000 ;
      LAYER met4 ;
        RECT 0.000000 29.500000 1.270000 34.150000 ;
      LAYER met5 ;
        RECT  25.935000 0.000000  30.385000 1.270000 ;
        RECT 175.785000 0.000000 200.000000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000  29.600000 1.270000  34.050000 ;
        RECT 0.000000 179.450000 1.270000 203.665000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 61.900000 1.270000 66.350000 ;
      LAYER met4 ;
        RECT 58.235000 0.000000 62.685000 1.270000 ;
      LAYER met5 ;
        RECT  0.000000 62.000000  1.270000 66.250000 ;
        RECT 58.335000  0.000000 62.585000  1.270000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 35.550000 1.270000 39.000000 ;
      LAYER met4 ;
        RECT 31.885000 0.000000 35.335000 1.270000 ;
      LAYER met5 ;
        RECT 0.000000 35.650000 1.270000 38.900000 ;
      LAYER met5 ;
        RECT 31.985000 0.000000 35.235000 1.270000 ;
    END
  END VSWITCH
END sky130_fd_io__corner_bus_overlay
END LIBRARY
