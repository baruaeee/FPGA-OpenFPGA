* NGSPICE file created from sky130_ef_sc_hd__newfill_12.ext - technology: sky130A

.subckt sky130_ef_sc_hd__newfill_12 VGND VPWR VPB VNB
.ends

