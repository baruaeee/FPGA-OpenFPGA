magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 3 21 735 203
rect 28 -17 62 21
<< scnmos >>
rect 81 47 111 177
rect 236 47 266 177
rect 338 47 368 177
rect 452 47 482 177
rect 555 47 585 177
rect 627 47 657 177
<< scpmoshvt >>
rect 81 297 111 497
rect 236 297 266 497
rect 338 297 368 497
rect 452 297 482 497
rect 537 297 567 497
rect 627 297 657 497
<< ndiff >>
rect 29 133 81 177
rect 29 99 37 133
rect 71 99 81 133
rect 29 47 81 99
rect 111 157 236 177
rect 111 55 121 157
rect 223 55 236 157
rect 111 47 236 55
rect 266 129 338 177
rect 266 95 285 129
rect 319 95 338 129
rect 266 47 338 95
rect 368 89 452 177
rect 368 55 393 89
rect 427 55 452 89
rect 368 47 452 55
rect 482 165 555 177
rect 482 131 502 165
rect 536 131 555 165
rect 482 97 555 131
rect 482 63 502 97
rect 536 63 555 97
rect 482 47 555 63
rect 585 47 627 177
rect 657 165 709 177
rect 657 131 667 165
rect 701 131 709 165
rect 657 97 709 131
rect 657 63 667 97
rect 701 63 709 97
rect 657 47 709 63
<< pdiff >>
rect 29 485 81 497
rect 29 451 37 485
rect 71 451 81 485
rect 29 417 81 451
rect 29 383 37 417
rect 71 383 81 417
rect 29 349 81 383
rect 29 315 37 349
rect 71 315 81 349
rect 29 297 81 315
rect 111 489 236 497
rect 111 455 148 489
rect 182 455 236 489
rect 111 421 236 455
rect 111 387 148 421
rect 182 387 236 421
rect 111 297 236 387
rect 266 297 338 497
rect 368 297 452 497
rect 482 489 537 497
rect 482 455 493 489
rect 527 455 537 489
rect 482 421 537 455
rect 482 387 493 421
rect 527 387 537 421
rect 482 353 537 387
rect 482 319 493 353
rect 527 319 537 353
rect 482 297 537 319
rect 567 485 627 497
rect 567 451 580 485
rect 614 451 627 485
rect 567 417 627 451
rect 567 383 580 417
rect 614 383 627 417
rect 567 297 627 383
rect 657 448 709 497
rect 657 414 667 448
rect 701 414 709 448
rect 657 380 709 414
rect 657 346 667 380
rect 701 346 709 380
rect 657 297 709 346
<< ndiffc >>
rect 37 99 71 133
rect 121 55 223 157
rect 285 95 319 129
rect 393 55 427 89
rect 502 131 536 165
rect 502 63 536 97
rect 667 131 701 165
rect 667 63 701 97
<< pdiffc >>
rect 37 451 71 485
rect 37 383 71 417
rect 37 315 71 349
rect 148 455 182 489
rect 148 387 182 421
rect 493 455 527 489
rect 493 387 527 421
rect 493 319 527 353
rect 580 451 614 485
rect 580 383 614 417
rect 667 414 701 448
rect 667 346 701 380
<< poly >>
rect 81 497 111 523
rect 236 497 266 523
rect 338 497 368 523
rect 452 497 482 523
rect 537 497 567 523
rect 627 497 657 523
rect 81 265 111 297
rect 236 265 266 297
rect 338 265 368 297
rect 452 265 482 297
rect 537 265 567 297
rect 627 265 657 297
rect 81 249 165 265
rect 81 215 121 249
rect 155 215 165 249
rect 81 199 165 215
rect 212 249 266 265
rect 212 215 222 249
rect 256 215 266 249
rect 212 199 266 215
rect 314 249 368 265
rect 314 215 324 249
rect 358 215 368 249
rect 314 199 368 215
rect 410 249 482 265
rect 410 215 420 249
rect 454 215 482 249
rect 410 199 482 215
rect 524 249 585 265
rect 524 215 534 249
rect 568 215 585 249
rect 524 199 585 215
rect 81 177 111 199
rect 236 177 266 199
rect 338 177 368 199
rect 452 177 482 199
rect 555 177 585 199
rect 627 249 715 265
rect 627 215 670 249
rect 704 215 715 249
rect 627 199 715 215
rect 627 177 657 199
rect 81 21 111 47
rect 236 21 266 47
rect 338 21 368 47
rect 452 21 482 47
rect 555 21 585 47
rect 627 21 657 47
<< polycont >>
rect 121 215 155 249
rect 222 215 256 249
rect 324 215 358 249
rect 420 215 454 249
rect 534 215 568 249
rect 670 215 704 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 485 87 493
rect 17 451 37 485
rect 71 451 87 485
rect 17 417 87 451
rect 17 383 37 417
rect 71 383 87 417
rect 17 349 87 383
rect 121 489 202 527
rect 121 455 148 489
rect 182 455 202 489
rect 121 421 202 455
rect 121 387 148 421
rect 182 387 202 421
rect 121 367 202 387
rect 236 489 543 493
rect 236 459 493 489
rect 17 315 37 349
rect 71 315 87 349
rect 236 333 270 459
rect 477 455 493 459
rect 527 455 543 489
rect 477 421 543 455
rect 17 214 87 315
rect 121 299 270 333
rect 121 249 155 299
rect 304 265 358 414
rect 17 133 71 214
rect 121 199 155 215
rect 189 249 256 265
rect 189 215 222 249
rect 189 199 256 215
rect 290 249 358 265
rect 290 215 324 249
rect 290 199 358 215
rect 396 265 443 414
rect 477 387 493 421
rect 527 387 543 421
rect 477 353 543 387
rect 580 485 627 527
rect 614 451 627 485
rect 580 417 627 451
rect 614 383 627 417
rect 580 367 627 383
rect 661 448 719 493
rect 661 414 667 448
rect 701 414 719 448
rect 661 380 719 414
rect 477 319 493 353
rect 527 333 543 353
rect 661 346 667 380
rect 701 346 719 380
rect 661 333 719 346
rect 527 319 719 333
rect 477 299 719 319
rect 396 249 454 265
rect 396 215 420 249
rect 396 199 454 215
rect 488 249 568 265
rect 488 215 534 249
rect 488 199 568 215
rect 602 165 636 299
rect 670 249 719 265
rect 704 215 719 249
rect 670 199 719 215
rect 17 99 37 133
rect 17 51 71 99
rect 105 157 239 165
rect 105 55 121 157
rect 223 55 239 157
rect 273 131 502 165
rect 536 131 552 165
rect 273 129 332 131
rect 273 95 285 129
rect 319 95 332 129
rect 486 97 552 131
rect 273 62 332 95
rect 368 89 443 97
rect 105 17 239 55
rect 368 55 393 89
rect 427 55 443 89
rect 486 63 502 97
rect 536 63 552 97
rect 486 62 552 63
rect 602 131 667 165
rect 701 131 719 165
rect 602 97 719 131
rect 602 63 667 97
rect 701 63 719 97
rect 368 17 443 55
rect 602 51 719 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 28 221 62 255 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 212 221 246 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 304 221 338 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 396 221 430 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 488 221 522 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 28 289 62 323 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 28 357 62 391 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 28 425 62 459 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 28 153 62 187 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 28 85 62 119 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 304 289 338 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 396 289 430 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 396 357 430 391 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 304 357 338 391 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o311a_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 920548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 912932
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 3.680 2.720 
<< end >>
