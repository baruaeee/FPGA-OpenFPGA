magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 551 203
rect 30 -17 64 21
<< locali >>
rect 19 459 253 493
rect 19 325 85 459
rect 187 451 253 459
rect 323 325 535 333
rect 19 299 535 325
rect 19 289 368 299
rect 25 153 115 255
rect 153 215 248 255
rect 198 135 248 215
rect 298 215 368 255
rect 298 135 340 215
rect 402 199 467 265
rect 501 165 535 299
rect 389 131 535 165
rect 389 101 425 131
rect 164 51 425 101
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 287 451 362 527
rect 119 417 165 425
rect 119 407 242 417
rect 391 407 425 433
rect 119 367 425 407
rect 472 371 525 527
rect 119 359 295 367
rect 19 17 109 119
rect 461 17 527 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 298 135 340 215 6 A1
port 1 nsew signal input
rlabel locali s 298 215 368 255 6 A1
port 1 nsew signal input
rlabel locali s 402 199 467 265 6 A2
port 2 nsew signal input
rlabel locali s 198 135 248 215 6 B1
port 3 nsew signal input
rlabel locali s 153 215 248 255 6 B1
port 3 nsew signal input
rlabel locali s 25 153 115 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 551 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 164 51 425 101 6 Y
port 9 nsew signal output
rlabel locali s 389 101 425 131 6 Y
port 9 nsew signal output
rlabel locali s 389 131 535 165 6 Y
port 9 nsew signal output
rlabel locali s 501 165 535 299 6 Y
port 9 nsew signal output
rlabel locali s 19 289 368 299 6 Y
port 9 nsew signal output
rlabel locali s 19 299 535 325 6 Y
port 9 nsew signal output
rlabel locali s 323 325 535 333 6 Y
port 9 nsew signal output
rlabel locali s 187 451 253 459 6 Y
port 9 nsew signal output
rlabel locali s 19 325 85 459 6 Y
port 9 nsew signal output
rlabel locali s 19 459 253 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4088784
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4083170
<< end >>
