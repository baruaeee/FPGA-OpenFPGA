magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 21 21 643 203
rect 29 -17 63 21
<< locali >>
rect 453 425 529 459
rect 495 391 529 425
rect 85 289 393 323
rect 85 199 134 289
rect 186 215 325 255
rect 359 249 393 289
rect 495 351 627 391
rect 359 215 479 249
rect 593 165 627 351
rect 563 69 627 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 425 77 527
rect 111 391 177 493
rect 211 425 337 527
rect 563 425 623 527
rect 17 357 461 391
rect 17 165 51 357
rect 427 317 461 357
rect 427 283 559 317
rect 525 199 559 283
rect 17 56 110 165
rect 211 17 245 181
rect 279 165 461 181
rect 279 147 529 165
rect 279 51 345 147
rect 427 131 529 147
rect 379 17 449 95
rect 483 51 529 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 186 215 325 255 6 A
port 1 nsew signal input
rlabel locali s 359 215 479 249 6 B
port 2 nsew signal input
rlabel locali s 359 249 393 289 6 B
port 2 nsew signal input
rlabel locali s 85 199 134 289 6 B
port 2 nsew signal input
rlabel locali s 85 289 393 323 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 21 21 643 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 563 69 627 165 6 Y
port 7 nsew signal output
rlabel locali s 593 165 627 351 6 Y
port 7 nsew signal output
rlabel locali s 495 351 627 391 6 Y
port 7 nsew signal output
rlabel locali s 495 391 529 425 6 Y
port 7 nsew signal output
rlabel locali s 453 425 529 459 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 624608
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 619304
<< end >>
