magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1365 157 1655 203
rect 1 21 1655 157
rect 29 -17 63 21
<< locali >>
rect 167 153 247 219
rect 204 79 247 153
rect 482 203 523 264
rect 448 143 523 203
rect 557 143 615 264
rect 949 143 1023 279
rect 1471 367 1553 491
rect 1491 299 1553 367
rect 1327 215 1389 265
rect 1307 199 1389 215
rect 1307 75 1369 199
rect 1519 145 1553 299
rect 1487 53 1553 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 35 417 69 475
rect 103 451 169 527
rect 282 425 448 459
rect 35 391 133 417
rect 35 383 380 391
rect 99 357 380 383
rect 29 323 65 349
rect 63 289 65 323
rect 29 195 65 289
rect 99 161 133 357
rect 201 289 213 323
rect 247 289 278 323
rect 244 257 278 289
rect 312 315 380 357
rect 34 127 133 161
rect 312 207 346 315
rect 414 281 448 425
rect 519 411 565 527
rect 661 425 764 459
rect 594 357 663 391
rect 713 362 764 425
rect 629 332 663 357
rect 629 298 683 332
rect 34 69 69 127
rect 103 17 169 93
rect 281 141 346 207
rect 380 247 448 281
rect 649 278 683 298
rect 380 107 414 247
rect 649 212 696 278
rect 294 73 414 107
rect 490 17 556 109
rect 649 93 683 212
rect 730 135 764 362
rect 597 59 683 93
rect 717 69 764 135
rect 798 425 903 459
rect 798 69 836 425
rect 951 401 1020 527
rect 1065 431 1255 465
rect 879 347 917 379
rect 1065 347 1099 431
rect 1305 425 1369 459
rect 879 313 1099 347
rect 879 117 913 313
rect 879 51 920 117
rect 959 17 1025 109
rect 1065 93 1099 313
rect 1133 207 1191 397
rect 1335 333 1369 425
rect 1403 367 1437 527
rect 1225 323 1293 329
rect 1259 289 1293 323
rect 1335 299 1457 333
rect 1587 299 1637 527
rect 1225 249 1293 289
rect 1423 265 1457 299
rect 1133 141 1257 207
rect 1423 199 1485 265
rect 1065 59 1244 93
rect 1403 17 1453 163
rect 1587 17 1638 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 289 63 323
rect 213 289 247 323
rect 1225 289 1259 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 17 323 75 329
rect 17 289 29 323
rect 63 320 75 323
rect 201 323 259 329
rect 201 320 213 323
rect 63 292 213 320
rect 63 289 75 292
rect 17 283 75 289
rect 201 289 213 292
rect 247 320 259 323
rect 1213 323 1271 329
rect 1213 320 1225 323
rect 247 292 1225 320
rect 247 289 259 292
rect 201 283 259 289
rect 1213 289 1225 292
rect 1259 289 1271 323
rect 1213 283 1271 289
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< obsm1 >>
rect 385 456 443 465
rect 661 456 719 465
rect 385 428 719 456
rect 385 419 443 428
rect 661 419 719 428
rect 845 456 903 465
rect 1305 456 1363 465
rect 845 428 1363 456
rect 845 419 903 428
rect 1305 419 1363 428
rect 293 388 351 397
rect 1121 388 1179 397
rect 293 360 1179 388
rect 293 351 351 360
rect 1121 351 1179 360
<< labels >>
rlabel locali s 1307 75 1369 199 6 A0
port 1 nsew signal input
rlabel locali s 1307 199 1389 215 6 A0
port 1 nsew signal input
rlabel locali s 1327 215 1389 265 6 A0
port 1 nsew signal input
rlabel locali s 949 143 1023 279 6 A1
port 2 nsew signal input
rlabel locali s 204 79 247 153 6 A2
port 3 nsew signal input
rlabel locali s 167 153 247 219 6 A2
port 3 nsew signal input
rlabel locali s 448 143 523 203 6 A3
port 4 nsew signal input
rlabel locali s 482 203 523 264 6 A3
port 4 nsew signal input
rlabel metal1 s 1213 283 1271 292 6 S0
port 5 nsew signal input
rlabel metal1 s 201 283 259 292 6 S0
port 5 nsew signal input
rlabel metal1 s 17 283 75 292 6 S0
port 5 nsew signal input
rlabel metal1 s 17 292 1271 320 6 S0
port 5 nsew signal input
rlabel metal1 s 1213 320 1271 329 6 S0
port 5 nsew signal input
rlabel metal1 s 201 320 259 329 6 S0
port 5 nsew signal input
rlabel metal1 s 17 320 75 329 6 S0
port 5 nsew signal input
rlabel locali s 557 143 615 264 6 S1
port 6 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1 21 1655 157 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1365 157 1655 203 6 VNB
port 8 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 1487 53 1553 145 6 X
port 11 nsew signal output
rlabel locali s 1519 145 1553 299 6 X
port 11 nsew signal output
rlabel locali s 1491 299 1553 367 6 X
port 11 nsew signal output
rlabel locali s 1471 367 1553 491 6 X
port 11 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1656 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1784296
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1770058
<< end >>
