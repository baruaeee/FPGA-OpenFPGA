magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 229 185 419 203
rect 33 21 419 185
rect 33 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 115 75 145 159
rect 199 75 229 159
rect 307 47 337 177
<< scpmoshvt >>
rect 115 371 145 455
rect 199 371 229 455
rect 307 297 337 497
<< ndiff >>
rect 255 159 307 177
rect 59 121 115 159
rect 59 87 71 121
rect 105 87 115 121
rect 59 75 115 87
rect 145 75 199 159
rect 229 93 307 159
rect 229 75 263 93
rect 255 59 263 75
rect 297 59 307 93
rect 255 47 307 59
rect 337 93 393 177
rect 337 59 347 93
rect 381 59 393 93
rect 337 47 393 59
<< pdiff >>
rect 255 485 307 497
rect 255 455 263 485
rect 59 443 115 455
rect 59 409 71 443
rect 105 409 115 443
rect 59 371 115 409
rect 145 443 199 455
rect 145 409 155 443
rect 189 409 199 443
rect 145 371 199 409
rect 229 451 263 455
rect 297 451 307 485
rect 229 417 307 451
rect 229 383 263 417
rect 297 383 307 417
rect 229 371 307 383
rect 245 297 307 371
rect 337 485 432 497
rect 337 451 367 485
rect 401 451 432 485
rect 337 417 432 451
rect 337 383 367 417
rect 401 383 432 417
rect 337 297 432 383
<< ndiffc >>
rect 71 87 105 121
rect 263 59 297 93
rect 347 59 381 93
<< pdiffc >>
rect 71 409 105 443
rect 155 409 189 443
rect 263 451 297 485
rect 263 383 297 417
rect 367 451 401 485
rect 367 383 401 417
<< poly >>
rect 307 497 337 523
rect 115 455 145 481
rect 199 455 229 481
rect 115 265 145 371
rect 58 249 145 265
rect 58 215 74 249
rect 108 215 145 249
rect 58 199 145 215
rect 115 159 145 199
rect 199 265 229 371
rect 307 265 337 297
rect 199 249 265 265
rect 199 215 215 249
rect 249 215 265 249
rect 199 199 265 215
rect 307 249 373 265
rect 307 215 323 249
rect 357 215 373 249
rect 307 199 373 215
rect 199 159 229 199
rect 307 177 337 199
rect 115 49 145 75
rect 199 49 229 75
rect 307 21 337 47
<< polycont >>
rect 74 215 108 249
rect 215 215 249 249
rect 323 215 357 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 57 443 113 527
rect 247 485 313 527
rect 57 409 71 443
rect 105 409 113 443
rect 57 393 113 409
rect 147 443 207 459
rect 147 409 155 443
rect 189 409 207 443
rect 147 349 207 409
rect 247 451 263 485
rect 297 451 313 485
rect 247 417 313 451
rect 247 383 263 417
rect 297 383 313 417
rect 351 485 443 493
rect 351 451 367 485
rect 401 451 443 485
rect 351 417 443 451
rect 351 383 367 417
rect 401 383 443 417
rect 20 265 73 337
rect 147 315 335 349
rect 301 265 335 315
rect 20 249 155 265
rect 20 215 74 249
rect 108 215 155 249
rect 199 249 267 265
rect 199 215 215 249
rect 249 215 267 249
rect 301 249 359 265
rect 301 215 323 249
rect 357 215 359 249
rect 301 199 359 215
rect 301 181 335 199
rect 57 143 335 181
rect 57 121 123 143
rect 57 87 71 121
rect 105 87 123 121
rect 393 109 443 383
rect 57 71 123 87
rect 247 93 297 109
rect 247 59 263 93
rect 247 17 297 59
rect 331 93 443 109
rect 331 59 347 93
rect 381 59 443 93
rect 331 51 443 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 397 153 431 187 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 85 431 119 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 289 431 323 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 357 431 391 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 425 431 459 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 SLEEP_B
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 lpflow_inputiso0n_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 2357562
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2352700
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 11.500 13.600 
<< end >>
