//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Template for user-defined Verilog modules
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Nov  3 15:48:23 2024
//-------------------------------------------
// ----- Template Verilog module for sky130_osu_sc_18T_hs__inv_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__inv_1 -----
module sky130_osu_sc_18T_hs__inv_1(A,
                                   Y);
//----- INPUT PORTS -----
input [0:0] A;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__inv_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_osu_sc_18T_hs__buf_4 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__buf_4 -----
module sky130_osu_sc_18T_hs__buf_4(A,
                                   Y);
//----- INPUT PORTS -----
input [0:0] A;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__buf_4 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_osu_sc_18T_hs__inv_4 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__inv_4 -----
module sky130_osu_sc_18T_hs__inv_4(A,
                                   Y);
//----- INPUT PORTS -----
input [0:0] A;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__inv_4 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_osu_sc_18T_hs__or2_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__or2_1 -----
module sky130_osu_sc_18T_hs__or2_1(A,
                                   B,
                                   Y);
//----- INPUT PORTS -----
input [0:0] A;
//----- INPUT PORTS -----
input [0:0] B;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__or2_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_osu_sc_18T_hs__mux2_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__mux2_1 -----
module sky130_osu_sc_18T_hs__mux2_1(A1,
                                    A0,
                                    S0,
                                    Y);
//----- INPUT PORTS -----
input [0:0] A1;
//----- INPUT PORTS -----
input [0:0] A0;
//----- INPUT PORTS -----
input [0:0] S0;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__mux2_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_osu_sc_18T_hs__dffsr_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__dffsr_1 -----
module sky130_osu_sc_18T_hs__dffsr_1(SN,
                                     RN,
                                     CK,
                                     D,
                                     Q);
//----- GLOBAL PORTS -----
input [0:0] SN;
//----- GLOBAL PORTS -----
input [0:0] RN;
//----- GLOBAL PORTS -----
input [0:0] CK;
//----- INPUT PORTS -----
input [0:0] D;
//----- OUTPUT PORTS -----
output [0:0] Q;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__dffsr_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_osu_sc_18T_hs__dffr_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_osu_sc_18T_hs__dffr_1 -----
module sky130_osu_sc_18T_hs__dffr_1(RN,
                                    CK,
                                    D,
                                    Q,
                                    QN);
//----- GLOBAL PORTS -----
input [0:0] RN;
//----- GLOBAL PORTS -----
input [0:0] CK;
//----- INPUT PORTS -----
input [0:0] D;
//----- OUTPUT PORTS -----
output [0:0] Q;
//----- OUTPUT PORTS -----
output [0:0] QN;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_osu_sc_18T_hs__dffr_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for GPIO -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for GPIO -----
module GPIO(PAD,
            A,
            DIR,
            Y);
//----- GPIO PORTS -----
inout [0:0] PAD;
//----- INPUT PORTS -----
input [0:0] A;
//----- INPUT PORTS -----
input [0:0] DIR;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for GPIO -----

//----- Default net type -----
`default_nettype wire


