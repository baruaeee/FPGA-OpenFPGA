/home/exotic/Desktop/FPGA-OpenFPGA/PNR/auto_3x3_sky_scl/lef/IO/sky130_fd_io__top_gpio_ovtv2.lef