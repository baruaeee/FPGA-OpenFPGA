magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1906 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1196 47 1226 177
rect 1280 47 1310 177
rect 1368 47 1398 177
rect 1452 47 1482 177
rect 1541 47 1571 177
rect 1625 47 1655 177
rect 1709 47 1739 177
rect 1793 47 1823 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 792 297 822 497
rect 876 297 906 497
rect 960 297 990 497
rect 1044 297 1074 497
rect 1133 297 1163 497
rect 1217 297 1247 497
rect 1301 297 1331 497
rect 1385 297 1415 497
rect 1571 297 1601 497
rect 1655 297 1685 497
rect 1739 297 1769 497
rect 1823 297 1853 497
<< ndiff >>
rect 27 95 79 177
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 47 163 129
rect 193 95 247 177
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 163 331 177
rect 277 129 287 163
rect 321 129 331 163
rect 277 47 331 129
rect 361 129 415 177
rect 361 95 371 129
rect 405 95 415 129
rect 361 47 415 95
rect 445 89 499 177
rect 445 55 455 89
rect 489 55 499 89
rect 445 47 499 55
rect 529 157 583 177
rect 529 123 539 157
rect 573 123 583 157
rect 529 47 583 123
rect 613 89 667 177
rect 613 55 623 89
rect 657 55 667 89
rect 613 47 667 55
rect 697 157 749 177
rect 697 123 707 157
rect 741 123 749 157
rect 697 47 749 123
rect 803 165 855 177
rect 803 131 811 165
rect 845 131 855 165
rect 803 47 855 131
rect 885 89 939 177
rect 885 55 895 89
rect 929 55 939 89
rect 885 47 939 55
rect 969 165 1023 177
rect 969 131 979 165
rect 1013 131 1023 165
rect 969 47 1023 131
rect 1053 89 1107 177
rect 1053 55 1063 89
rect 1097 55 1107 89
rect 1053 47 1107 55
rect 1137 165 1196 177
rect 1137 131 1152 165
rect 1186 131 1196 165
rect 1137 47 1196 131
rect 1226 93 1280 177
rect 1226 59 1236 93
rect 1270 59 1280 93
rect 1226 47 1280 59
rect 1310 165 1368 177
rect 1310 131 1320 165
rect 1354 131 1368 165
rect 1310 47 1368 131
rect 1398 90 1452 177
rect 1398 56 1408 90
rect 1442 56 1452 90
rect 1398 47 1452 56
rect 1482 165 1541 177
rect 1482 131 1497 165
rect 1531 131 1541 165
rect 1482 47 1541 131
rect 1571 89 1625 177
rect 1571 55 1581 89
rect 1615 55 1625 89
rect 1571 47 1625 55
rect 1655 165 1709 177
rect 1655 131 1665 165
rect 1699 131 1709 165
rect 1655 47 1709 131
rect 1739 89 1793 177
rect 1739 55 1749 89
rect 1783 55 1793 89
rect 1739 47 1793 55
rect 1823 165 1880 177
rect 1823 131 1833 165
rect 1867 131 1880 165
rect 1823 47 1880 131
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 421 163 455
rect 109 387 119 421
rect 153 387 163 421
rect 109 297 163 387
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 489 331 497
rect 277 455 287 489
rect 321 455 331 489
rect 277 421 331 455
rect 277 387 287 421
rect 321 387 331 421
rect 277 297 331 387
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 489 499 497
rect 445 455 455 489
rect 489 455 499 489
rect 445 421 499 455
rect 445 387 455 421
rect 489 387 499 421
rect 445 297 499 387
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 409 583 443
rect 529 375 539 409
rect 573 375 583 409
rect 529 297 583 375
rect 613 489 667 497
rect 613 455 623 489
rect 657 455 667 489
rect 613 421 667 455
rect 613 387 623 421
rect 657 387 667 421
rect 613 297 667 387
rect 697 477 792 497
rect 697 443 707 477
rect 741 443 792 477
rect 697 409 792 443
rect 697 375 707 409
rect 741 375 792 409
rect 697 297 792 375
rect 822 489 876 497
rect 822 455 832 489
rect 866 455 876 489
rect 822 421 876 455
rect 822 387 832 421
rect 866 387 876 421
rect 822 297 876 387
rect 906 477 960 497
rect 906 443 916 477
rect 950 443 960 477
rect 906 409 960 443
rect 906 375 916 409
rect 950 375 960 409
rect 906 297 960 375
rect 990 489 1044 497
rect 990 455 1000 489
rect 1034 455 1044 489
rect 990 421 1044 455
rect 990 387 1000 421
rect 1034 387 1044 421
rect 990 297 1044 387
rect 1074 477 1133 497
rect 1074 443 1084 477
rect 1118 443 1133 477
rect 1074 409 1133 443
rect 1074 375 1084 409
rect 1118 375 1133 409
rect 1074 297 1133 375
rect 1163 489 1217 497
rect 1163 455 1173 489
rect 1207 455 1217 489
rect 1163 421 1217 455
rect 1163 387 1173 421
rect 1207 387 1217 421
rect 1163 297 1217 387
rect 1247 404 1301 497
rect 1247 370 1257 404
rect 1291 370 1301 404
rect 1247 297 1301 370
rect 1331 443 1385 497
rect 1331 409 1341 443
rect 1375 409 1385 443
rect 1331 297 1385 409
rect 1415 364 1465 497
rect 1519 485 1571 497
rect 1519 451 1527 485
rect 1561 451 1571 485
rect 1519 440 1571 451
rect 1415 343 1467 364
rect 1415 309 1425 343
rect 1459 309 1467 343
rect 1415 297 1467 309
rect 1521 297 1571 440
rect 1601 477 1655 497
rect 1601 443 1611 477
rect 1645 443 1655 477
rect 1601 409 1655 443
rect 1601 375 1611 409
rect 1645 375 1655 409
rect 1601 297 1655 375
rect 1685 489 1739 497
rect 1685 455 1695 489
rect 1729 455 1739 489
rect 1685 421 1739 455
rect 1685 387 1695 421
rect 1729 387 1739 421
rect 1685 297 1739 387
rect 1769 477 1823 497
rect 1769 443 1779 477
rect 1813 443 1823 477
rect 1769 409 1823 443
rect 1769 375 1779 409
rect 1813 375 1823 409
rect 1769 297 1823 375
rect 1853 485 1905 497
rect 1853 451 1863 485
rect 1897 451 1905 485
rect 1853 417 1905 451
rect 1853 383 1863 417
rect 1897 383 1905 417
rect 1853 297 1905 383
<< ndiffc >>
rect 35 61 69 95
rect 119 129 153 163
rect 203 61 237 95
rect 287 129 321 163
rect 371 95 405 129
rect 455 55 489 89
rect 539 123 573 157
rect 623 55 657 89
rect 707 123 741 157
rect 811 131 845 165
rect 895 55 929 89
rect 979 131 1013 165
rect 1063 55 1097 89
rect 1152 131 1186 165
rect 1236 59 1270 93
rect 1320 131 1354 165
rect 1408 56 1442 90
rect 1497 131 1531 165
rect 1581 55 1615 89
rect 1665 131 1699 165
rect 1749 55 1783 89
rect 1833 131 1867 165
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 455 153 489
rect 119 387 153 421
rect 203 443 237 477
rect 203 375 237 409
rect 287 455 321 489
rect 287 387 321 421
rect 371 443 405 477
rect 371 375 405 409
rect 455 455 489 489
rect 455 387 489 421
rect 539 443 573 477
rect 539 375 573 409
rect 623 455 657 489
rect 623 387 657 421
rect 707 443 741 477
rect 707 375 741 409
rect 832 455 866 489
rect 832 387 866 421
rect 916 443 950 477
rect 916 375 950 409
rect 1000 455 1034 489
rect 1000 387 1034 421
rect 1084 443 1118 477
rect 1084 375 1118 409
rect 1173 455 1207 489
rect 1173 387 1207 421
rect 1257 370 1291 404
rect 1341 409 1375 443
rect 1527 451 1561 485
rect 1425 309 1459 343
rect 1611 443 1645 477
rect 1611 375 1645 409
rect 1695 455 1729 489
rect 1695 387 1729 421
rect 1779 443 1813 477
rect 1779 375 1813 409
rect 1863 451 1897 485
rect 1863 383 1897 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 792 497 822 523
rect 876 497 906 523
rect 960 497 990 523
rect 1044 497 1074 523
rect 1133 497 1163 523
rect 1217 497 1247 523
rect 1301 497 1331 523
rect 1385 497 1415 523
rect 1571 497 1601 523
rect 1655 497 1685 523
rect 1739 497 1769 523
rect 1823 497 1853 523
rect 79 277 109 297
rect 163 277 193 297
rect 247 277 277 297
rect 331 277 361 297
rect 79 249 361 277
rect 79 215 125 249
rect 159 215 207 249
rect 241 215 296 249
rect 330 215 361 249
rect 79 205 361 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 792 259 822 297
rect 876 259 906 297
rect 960 259 990 297
rect 1044 259 1074 297
rect 1133 282 1163 297
rect 1217 282 1247 297
rect 1133 263 1247 282
rect 1139 262 1247 263
rect 1140 261 1247 262
rect 1141 260 1247 261
rect 1142 259 1247 260
rect 1301 259 1331 297
rect 1385 259 1415 297
rect 1571 259 1601 297
rect 1655 259 1685 297
rect 1739 259 1769 297
rect 1823 259 1853 297
rect 415 249 697 259
rect 415 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 697 249
rect 415 205 697 215
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 776 249 1074 259
rect 1143 258 1482 259
rect 1145 257 1482 258
rect 1146 256 1482 257
rect 1148 255 1482 256
rect 1149 254 1482 255
rect 1152 253 1482 254
rect 1155 252 1482 253
rect 776 215 834 249
rect 868 215 902 249
rect 936 215 970 249
rect 1004 222 1074 249
rect 1196 249 1482 252
rect 1004 221 1115 222
rect 1004 220 1118 221
rect 1004 219 1121 220
rect 1004 218 1122 219
rect 1004 217 1124 218
rect 1004 216 1125 217
rect 1004 215 1127 216
rect 1196 215 1246 249
rect 1280 215 1314 249
rect 1348 215 1382 249
rect 1416 215 1482 249
rect 776 214 1128 215
rect 776 213 1129 214
rect 776 204 1137 213
rect 855 177 885 204
rect 939 177 969 204
rect 1023 192 1137 204
rect 1023 177 1053 192
rect 1107 177 1137 192
rect 1196 205 1482 215
rect 1196 177 1226 205
rect 1280 177 1310 205
rect 1368 177 1398 205
rect 1452 177 1482 205
rect 1541 249 1854 259
rect 1541 215 1581 249
rect 1615 215 1649 249
rect 1683 215 1717 249
rect 1751 215 1785 249
rect 1819 215 1854 249
rect 1541 205 1854 215
rect 1541 177 1571 205
rect 1625 177 1655 205
rect 1709 177 1739 205
rect 1793 177 1823 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1196 21 1226 47
rect 1280 21 1310 47
rect 1368 21 1398 47
rect 1452 21 1482 47
rect 1541 21 1571 47
rect 1625 21 1655 47
rect 1709 21 1739 47
rect 1793 21 1823 47
<< polycont >>
rect 125 215 159 249
rect 207 215 241 249
rect 296 215 330 249
rect 431 215 465 249
rect 499 215 533 249
rect 567 215 601 249
rect 635 215 669 249
rect 834 215 868 249
rect 902 215 936 249
rect 970 215 1004 249
rect 1246 215 1280 249
rect 1314 215 1348 249
rect 1382 215 1416 249
rect 1581 215 1615 249
rect 1649 215 1683 249
rect 1717 215 1751 249
rect 1785 215 1819 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 477 72 493
rect 17 443 35 477
rect 69 443 72 477
rect 17 409 72 443
rect 17 375 35 409
rect 69 375 72 409
rect 17 337 72 375
rect 106 489 169 527
rect 106 455 119 489
rect 153 455 169 489
rect 106 421 169 455
rect 106 387 119 421
rect 153 387 169 421
rect 106 371 169 387
rect 203 477 239 493
rect 237 443 239 477
rect 203 409 239 443
rect 237 375 239 409
rect 203 337 239 375
rect 278 489 335 527
rect 278 455 287 489
rect 321 455 335 489
rect 278 421 335 455
rect 278 387 287 421
rect 321 387 335 421
rect 278 371 335 387
rect 369 477 407 493
rect 369 443 371 477
rect 405 443 407 477
rect 369 409 407 443
rect 369 375 371 409
rect 405 375 407 409
rect 369 337 407 375
rect 441 489 503 527
rect 441 455 455 489
rect 489 455 503 489
rect 441 421 503 455
rect 441 387 455 421
rect 489 387 503 421
rect 441 371 503 387
rect 537 477 575 493
rect 537 443 539 477
rect 573 443 575 477
rect 537 409 575 443
rect 537 375 539 409
rect 573 375 575 409
rect 537 337 575 375
rect 609 489 671 527
rect 609 455 623 489
rect 657 455 671 489
rect 609 421 671 455
rect 609 387 623 421
rect 657 387 671 421
rect 609 371 671 387
rect 705 477 743 493
rect 705 443 707 477
rect 741 443 743 477
rect 705 409 743 443
rect 705 375 707 409
rect 741 375 743 409
rect 705 337 743 375
rect 815 489 880 527
rect 815 455 832 489
rect 866 455 880 489
rect 815 421 880 455
rect 815 387 832 421
rect 866 387 880 421
rect 815 371 880 387
rect 914 477 952 493
rect 914 443 916 477
rect 950 443 952 477
rect 914 409 952 443
rect 914 375 916 409
rect 950 375 952 409
rect 914 337 952 375
rect 986 489 1044 527
rect 986 455 1000 489
rect 1034 455 1044 489
rect 986 421 1044 455
rect 986 387 1000 421
rect 1034 387 1044 421
rect 986 371 1044 387
rect 1082 477 1120 493
rect 1082 443 1084 477
rect 1118 443 1120 477
rect 1082 409 1120 443
rect 1082 375 1084 409
rect 1118 375 1120 409
rect 1082 337 1120 375
rect 1157 489 1401 493
rect 1157 455 1173 489
rect 1207 455 1401 489
rect 1157 454 1401 455
rect 1157 421 1223 454
rect 1157 387 1173 421
rect 1207 387 1223 421
rect 1341 443 1401 454
rect 1511 485 1577 527
rect 1511 451 1527 485
rect 1561 451 1577 485
rect 1511 446 1577 451
rect 1611 477 1647 493
rect 1157 371 1223 387
rect 1257 404 1296 420
rect 1291 370 1296 404
rect 1375 412 1401 443
rect 1645 443 1647 477
rect 1611 412 1647 443
rect 1375 409 1647 412
rect 1341 378 1611 409
rect 1257 337 1296 370
rect 1609 375 1611 378
rect 1645 375 1647 409
rect 1409 343 1478 344
rect 1409 337 1425 343
rect 17 309 1425 337
rect 1459 309 1478 343
rect 17 303 1478 309
rect 1609 337 1647 375
rect 1682 489 1744 527
rect 1682 455 1695 489
rect 1729 455 1744 489
rect 1682 421 1744 455
rect 1682 387 1695 421
rect 1729 387 1744 421
rect 1682 371 1744 387
rect 1778 477 1816 493
rect 1778 443 1779 477
rect 1813 443 1816 477
rect 1778 409 1816 443
rect 1778 375 1779 409
rect 1813 375 1816 409
rect 1778 337 1816 375
rect 1609 303 1816 337
rect 1853 485 1915 527
rect 1853 451 1863 485
rect 1897 451 1915 485
rect 1853 417 1915 451
rect 1853 383 1863 417
rect 1897 383 1915 417
rect 1853 307 1915 383
rect 17 163 75 303
rect 109 249 351 269
rect 109 215 125 249
rect 159 215 207 249
rect 241 215 296 249
rect 330 215 351 249
rect 388 249 710 269
rect 388 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 710 249
rect 763 249 1091 269
rect 763 215 834 249
rect 868 215 902 249
rect 936 215 970 249
rect 1004 215 1091 249
rect 1222 249 1465 269
rect 1222 215 1246 249
rect 1280 215 1314 249
rect 1348 215 1382 249
rect 1416 215 1465 249
rect 1564 249 1915 268
rect 1564 215 1581 249
rect 1615 215 1649 249
rect 1683 215 1717 249
rect 1751 215 1785 249
rect 1819 215 1915 249
rect 795 165 1888 181
rect 17 129 119 163
rect 153 129 287 163
rect 321 129 337 163
rect 371 157 757 165
rect 371 129 539 157
rect 405 123 539 129
rect 573 123 707 157
rect 741 123 757 157
rect 795 131 811 165
rect 845 131 979 165
rect 1013 131 1152 165
rect 1186 131 1320 165
rect 1354 131 1497 165
rect 1531 131 1665 165
rect 1699 131 1833 165
rect 1867 131 1888 165
rect 19 61 35 95
rect 69 61 203 95
rect 237 61 405 95
rect 1220 93 1286 97
rect 19 57 405 61
rect 439 55 455 89
rect 489 55 623 89
rect 657 55 895 89
rect 929 55 1063 89
rect 1097 55 1113 89
rect 439 51 1113 55
rect 1220 59 1236 93
rect 1270 59 1286 93
rect 1220 17 1286 59
rect 1392 90 1458 97
rect 1392 56 1408 90
rect 1442 56 1458 90
rect 1392 17 1458 56
rect 1565 89 1631 97
rect 1565 55 1581 89
rect 1615 55 1631 89
rect 1565 17 1631 55
rect 1733 89 1799 97
rect 1733 55 1749 89
rect 1783 55 1799 89
rect 1733 17 1799 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 1869 221 1903 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 1777 221 1811 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 1685 221 1719 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 1593 221 1627 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 1409 221 1443 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 153 64 187 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 30 425 64 459 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o2111ai_4
rlabel metal1 s 0 -48 1932 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 976088
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 960678
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 9.660 2.720 
<< end >>
