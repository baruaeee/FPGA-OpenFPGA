/home/cae1/Desktop/FPGA-OpenFPGA/PNR/auto_3x3/lef/sky130_fd_sc_hd.lef