magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 544 157 827 203
rect 21 21 827 157
rect 29 -17 63 21
<< scnmos >>
rect 99 47 129 131
rect 171 47 201 131
rect 255 47 285 131
rect 327 47 357 131
rect 411 47 441 131
rect 483 47 513 131
rect 633 47 663 177
rect 717 47 747 177
<< scpmoshvt >>
rect 99 369 129 497
rect 171 369 201 497
rect 255 369 285 497
rect 327 369 357 497
rect 411 369 441 497
rect 483 369 513 497
rect 633 297 663 497
rect 717 297 747 497
<< ndiff >>
rect 570 131 633 177
rect 47 106 99 131
rect 47 72 55 106
rect 89 72 99 106
rect 47 47 99 72
rect 129 47 171 131
rect 201 89 255 131
rect 201 55 211 89
rect 245 55 255 89
rect 201 47 255 55
rect 285 47 327 131
rect 357 89 411 131
rect 357 55 367 89
rect 401 55 411 89
rect 357 47 411 55
rect 441 47 483 131
rect 513 93 633 131
rect 513 59 543 93
rect 577 59 633 93
rect 513 47 633 59
rect 663 165 717 177
rect 663 131 673 165
rect 707 131 717 165
rect 663 97 717 131
rect 663 63 673 97
rect 707 63 717 97
rect 663 47 717 63
rect 747 165 801 177
rect 747 131 757 165
rect 791 131 801 165
rect 747 97 801 131
rect 747 63 757 97
rect 791 63 801 97
rect 747 47 801 63
<< pdiff >>
rect 47 485 99 497
rect 47 451 55 485
rect 89 451 99 485
rect 47 417 99 451
rect 47 383 55 417
rect 89 383 99 417
rect 47 369 99 383
rect 129 369 171 497
rect 201 485 255 497
rect 201 451 211 485
rect 245 451 255 485
rect 201 369 255 451
rect 285 369 327 497
rect 357 485 411 497
rect 357 451 367 485
rect 401 451 411 485
rect 357 417 411 451
rect 357 383 367 417
rect 401 383 411 417
rect 357 369 411 383
rect 441 369 483 497
rect 513 485 633 497
rect 513 451 523 485
rect 557 451 633 485
rect 513 417 633 451
rect 513 383 523 417
rect 557 383 633 417
rect 513 369 633 383
rect 583 297 633 369
rect 663 485 717 497
rect 663 451 673 485
rect 707 451 717 485
rect 663 417 717 451
rect 663 383 673 417
rect 707 383 717 417
rect 663 349 717 383
rect 663 315 673 349
rect 707 315 717 349
rect 663 297 717 315
rect 747 485 801 497
rect 747 451 757 485
rect 791 451 801 485
rect 747 417 801 451
rect 747 383 757 417
rect 791 383 801 417
rect 747 349 801 383
rect 747 315 757 349
rect 791 315 801 349
rect 747 297 801 315
<< ndiffc >>
rect 55 72 89 106
rect 211 55 245 89
rect 367 55 401 89
rect 543 59 577 93
rect 673 131 707 165
rect 673 63 707 97
rect 757 131 791 165
rect 757 63 791 97
<< pdiffc >>
rect 55 451 89 485
rect 55 383 89 417
rect 211 451 245 485
rect 367 451 401 485
rect 367 383 401 417
rect 523 451 557 485
rect 523 383 557 417
rect 673 451 707 485
rect 673 383 707 417
rect 673 315 707 349
rect 757 451 791 485
rect 757 383 791 417
rect 757 315 791 349
<< poly >>
rect 99 497 129 523
rect 171 497 201 523
rect 255 497 285 523
rect 327 497 357 523
rect 411 497 441 523
rect 483 497 513 523
rect 633 497 663 523
rect 717 497 747 523
rect 99 265 129 369
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 99 131 129 199
rect 171 265 201 369
rect 255 265 285 369
rect 171 249 285 265
rect 171 215 211 249
rect 245 215 285 249
rect 171 199 285 215
rect 171 131 201 199
rect 255 131 285 199
rect 327 265 357 369
rect 411 265 441 369
rect 327 249 441 265
rect 327 215 373 249
rect 407 215 441 249
rect 327 199 441 215
rect 327 131 357 199
rect 411 131 441 199
rect 483 331 513 369
rect 483 321 549 331
rect 483 287 499 321
rect 533 287 549 321
rect 483 277 549 287
rect 483 131 513 277
rect 633 259 663 297
rect 717 259 747 297
rect 589 249 747 259
rect 589 215 605 249
rect 639 215 747 249
rect 589 205 747 215
rect 633 177 663 205
rect 717 177 747 205
rect 99 21 129 47
rect 171 21 201 47
rect 255 21 285 47
rect 327 21 357 47
rect 411 21 441 47
rect 483 21 513 47
rect 633 21 663 47
rect 717 21 747 47
<< polycont >>
rect 85 215 119 249
rect 211 215 245 249
rect 373 215 407 249
rect 499 287 533 321
rect 605 215 639 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 485 123 493
rect 17 451 55 485
rect 89 451 123 485
rect 17 417 123 451
rect 195 485 261 527
rect 195 451 211 485
rect 245 451 261 485
rect 195 435 261 451
rect 351 485 417 493
rect 351 451 367 485
rect 401 451 417 485
rect 17 383 55 417
rect 89 401 123 417
rect 351 417 417 451
rect 351 401 367 417
rect 89 383 367 401
rect 401 383 417 417
rect 17 367 417 383
rect 507 485 572 527
rect 507 451 523 485
rect 557 451 572 485
rect 507 417 572 451
rect 507 383 523 417
rect 557 383 572 417
rect 507 367 572 383
rect 657 485 723 493
rect 657 451 673 485
rect 707 451 723 485
rect 657 417 723 451
rect 657 383 673 417
rect 707 383 723 417
rect 17 165 51 367
rect 657 349 723 383
rect 85 321 614 333
rect 85 299 499 321
rect 85 249 155 299
rect 483 287 499 299
rect 533 287 614 321
rect 657 315 673 349
rect 707 315 723 349
rect 657 299 723 315
rect 757 485 811 527
rect 791 451 811 485
rect 757 417 811 451
rect 791 383 811 417
rect 757 349 811 383
rect 791 315 811 349
rect 757 299 811 315
rect 483 283 614 287
rect 119 215 155 249
rect 85 199 155 215
rect 201 249 339 265
rect 201 215 211 249
rect 245 215 339 249
rect 201 199 339 215
rect 373 249 431 265
rect 407 215 431 249
rect 373 199 431 215
rect 585 215 605 249
rect 639 215 655 249
rect 585 165 621 215
rect 689 181 723 299
rect 17 131 621 165
rect 657 165 723 181
rect 657 131 673 165
rect 707 131 723 165
rect 17 106 105 131
rect 17 72 55 106
rect 89 72 105 106
rect 17 56 105 72
rect 195 89 261 97
rect 195 55 211 89
rect 245 55 261 89
rect 195 17 261 55
rect 351 89 417 131
rect 657 97 723 131
rect 351 55 367 89
rect 401 55 417 89
rect 351 51 417 55
rect 527 93 593 97
rect 527 59 543 93
rect 577 59 593 93
rect 527 17 593 59
rect 657 63 673 97
rect 707 63 723 97
rect 657 51 723 63
rect 757 165 811 181
rect 791 131 811 165
rect 757 97 811 131
rect 791 63 811 97
rect 757 17 811 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 580 289 614 323 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 672 85 706 119 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
rlabel comment s 0 0 0 0 4 maj3_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1660154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1653706
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
