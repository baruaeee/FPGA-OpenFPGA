//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Template for user-defined Verilog modules
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat Oct 26 04:14:15 2024
//-------------------------------------------
// ----- Template Verilog module for sky130_fd_sc_hd__inv_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__inv_1 -----
module sky130_fd_sc_hd__inv_1(A,
                              Y);
//----- INPUT PORTS -----
input [0:0] A;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__inv_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_fd_sc_hd__buf_4 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__buf_4 -----
module sky130_fd_sc_hd__buf_4(A,
                              X);
//----- INPUT PORTS -----
input [0:0] A;
//----- OUTPUT PORTS -----
output [0:0] X;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__buf_4 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_fd_sc_hd__inv_4 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__inv_4 -----
module sky130_fd_sc_hd__inv_4(A,
                              Y);
//----- INPUT PORTS -----
input [0:0] A;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__inv_4 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_fd_sc_hd__or2_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__or2_1 -----
module sky130_fd_sc_hd__or2_1(A,
                              B,
                              X);
//----- INPUT PORTS -----
input [0:0] A;
//----- INPUT PORTS -----
input [0:0] B;
//----- OUTPUT PORTS -----
output [0:0] X;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__or2_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_fd_sc_hd__mux2_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__mux2_1 -----
module sky130_fd_sc_hd__mux2_1(A1,
                               A0,
                               S,
                               X);
//----- INPUT PORTS -----
input [0:0] A1;
//----- INPUT PORTS -----
input [0:0] A0;
//----- INPUT PORTS -----
input [0:0] S;
//----- OUTPUT PORTS -----
output [0:0] X;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__mux2_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_fd_sc_hd__sdfbbp_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__sdfbbp_1 -----
module sky130_fd_sc_hd__sdfbbp_1(SET_B,
                                 RESET_B,
                                 CLK,
                                 D,
                                 Q);
//----- GLOBAL PORTS -----
input [0:0] SET_B;
//----- GLOBAL PORTS -----
input [0:0] RESET_B;
//----- GLOBAL PORTS -----
input [0:0] CLK;
//----- INPUT PORTS -----
input [0:0] D;
//----- OUTPUT PORTS -----
output [0:0] Q;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__sdfbbp_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for sky130_fd_sc_hd__dfrbp_1 -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sky130_fd_sc_hd__dfrbp_1 -----
module sky130_fd_sc_hd__dfrbp_1(RESET_B,
                                CLK,
                                D,
                                Q,
                                Q_N);
//----- GLOBAL PORTS -----
input [0:0] RESET_B;
//----- GLOBAL PORTS -----
input [0:0] CLK;
//----- INPUT PORTS -----
input [0:0] D;
//----- OUTPUT PORTS -----
output [0:0] Q;
//----- OUTPUT PORTS -----
output [0:0] Q_N;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for sky130_fd_sc_hd__dfrbp_1 -----

//----- Default net type -----
`default_nettype wire


// ----- Template Verilog module for GPIO -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for GPIO -----
module GPIO(PAD,
            A,
            DIR,
            Y);
//----- GPIO PORTS -----
inout [0:0] PAD;
//----- INPUT PORTS -----
input [0:0] A;
//----- INPUT PORTS -----
input [0:0] DIR;
//----- OUTPUT PORTS -----
output [0:0] Y;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----

// ----- Internal logic should start here -----


// ----- Internal logic should end here -----
endmodule
// ----- END Verilog module for GPIO -----

//----- Default net type -----
`default_nettype wire


