/home/exotic/Desktop/FPGA-OpenFPGA/PNR/auto_3x3_gpdk/techlef/gsclib045_tech.lef