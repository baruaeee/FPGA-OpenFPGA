magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 7 21 1309 203
rect 29 -17 63 21
<< locali >>
rect 213 325 255 493
rect 373 325 423 493
rect 645 325 695 425
rect 813 325 863 425
rect 213 291 863 325
rect 489 289 863 291
rect 17 215 111 257
rect 489 215 579 289
rect 1317 257 1362 491
rect 613 215 895 255
rect 929 215 1362 257
rect 489 163 535 215
rect 284 129 535 163
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 29 325 95 487
rect 129 359 171 527
rect 289 359 339 527
rect 457 359 507 527
rect 555 459 947 493
rect 555 359 611 459
rect 729 359 779 459
rect 29 291 179 325
rect 897 325 947 459
rect 981 359 1031 527
rect 1065 325 1115 493
rect 1149 359 1199 527
rect 1233 325 1283 493
rect 897 291 1283 325
rect 145 257 179 291
rect 145 215 455 257
rect 145 179 179 215
rect 45 17 79 179
rect 113 58 179 179
rect 569 145 1291 181
rect 569 95 619 145
rect 216 61 619 95
rect 653 17 687 111
rect 721 51 787 145
rect 821 17 855 111
rect 889 51 955 145
rect 989 17 1023 111
rect 1057 51 1123 145
rect 1157 17 1191 111
rect 1225 51 1291 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
rlabel locali s 929 215 1362 257 6 A1
port 1 nsew signal input
rlabel locali s 1317 257 1362 491 6 A1
port 1 nsew signal input
rlabel locali s 613 215 895 255 6 A2
port 2 nsew signal input
rlabel locali s 17 215 111 257 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 7 21 1309 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 284 129 535 163 6 Y
port 8 nsew signal output
rlabel locali s 489 163 535 215 6 Y
port 8 nsew signal output
rlabel locali s 489 215 579 289 6 Y
port 8 nsew signal output
rlabel locali s 489 289 863 291 6 Y
port 8 nsew signal output
rlabel locali s 213 291 863 325 6 Y
port 8 nsew signal output
rlabel locali s 813 325 863 425 6 Y
port 8 nsew signal output
rlabel locali s 645 325 695 425 6 Y
port 8 nsew signal output
rlabel locali s 373 325 423 493 6 Y
port 8 nsew signal output
rlabel locali s 213 325 255 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1380 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1352826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1342018
<< end >>
