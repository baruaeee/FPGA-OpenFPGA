magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 157 604 203
rect 1 67 827 157
rect 29 21 827 67
rect 29 -17 63 21
<< locali >>
rect 224 333 290 493
rect 428 333 494 493
rect 86 215 156 331
rect 224 299 534 333
rect 194 215 264 265
rect 300 147 344 265
rect 484 165 534 299
rect 484 51 586 165
rect 678 145 728 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 413 85 493
rect 17 181 52 413
rect 119 367 185 527
rect 328 367 394 527
rect 536 435 690 527
rect 727 401 811 493
rect 568 367 811 401
rect 17 143 254 181
rect 17 97 85 143
rect 216 111 254 143
rect 394 111 450 265
rect 119 17 180 109
rect 216 73 450 111
rect 568 199 618 367
rect 762 109 811 367
rect 620 17 690 109
rect 724 51 811 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 678 145 728 323 6 A_N
port 1 nsew signal input
rlabel locali s 86 215 156 331 6 B_N
port 2 nsew signal input
rlabel locali s 300 147 344 265 6 C
port 3 nsew signal input
rlabel locali s 194 215 264 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 29 21 827 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 67 827 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 157 604 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 484 51 586 165 6 Y
port 9 nsew signal output
rlabel locali s 484 165 534 299 6 Y
port 9 nsew signal output
rlabel locali s 224 299 534 333 6 Y
port 9 nsew signal output
rlabel locali s 428 333 494 493 6 Y
port 9 nsew signal output
rlabel locali s 224 333 290 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1933288
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1926132
<< end >>
