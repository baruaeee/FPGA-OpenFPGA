magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 34 21 808 203
rect 34 17 63 21
rect 29 -17 63 17
<< locali >>
rect 136 333 202 493
rect 304 333 370 493
rect 472 333 538 493
rect 640 333 706 493
rect 17 299 811 333
rect 17 181 86 299
rect 136 215 707 265
rect 747 181 811 299
rect 17 143 811 181
rect 136 51 202 143
rect 304 51 370 143
rect 472 51 538 143
rect 640 51 706 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 51 367 102 527
rect 236 367 270 527
rect 404 367 438 527
rect 572 367 606 527
rect 740 367 800 527
rect 51 17 102 109
rect 236 17 270 109
rect 404 17 438 109
rect 572 17 606 109
rect 740 17 801 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 136 215 707 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 34 17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 34 21 808 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 640 51 706 143 6 Y
port 6 nsew signal output
rlabel locali s 472 51 538 143 6 Y
port 6 nsew signal output
rlabel locali s 304 51 370 143 6 Y
port 6 nsew signal output
rlabel locali s 136 51 202 143 6 Y
port 6 nsew signal output
rlabel locali s 17 143 811 181 6 Y
port 6 nsew signal output
rlabel locali s 747 181 811 299 6 Y
port 6 nsew signal output
rlabel locali s 17 181 86 299 6 Y
port 6 nsew signal output
rlabel locali s 17 299 811 333 6 Y
port 6 nsew signal output
rlabel locali s 640 333 706 493 6 Y
port 6 nsew signal output
rlabel locali s 472 333 538 493 6 Y
port 6 nsew signal output
rlabel locali s 304 333 370 493 6 Y
port 6 nsew signal output
rlabel locali s 136 333 202 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2208764
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2201264
<< end >>
