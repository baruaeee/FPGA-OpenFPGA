# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_gpio_ovtv2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 140 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  215.1680 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 53.125000 140.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  215.1680 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 48.365000 140.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    ANTENNAPARTIALCUTAREA  0.320000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.930000 14.070000 8.710000 14.390000 ;
        RECT 7.935000 14.065000 8.705000 14.070000 ;
        RECT 8.025000 13.975000 8.615000 14.065000 ;
        RECT 8.115000  0.000000 8.445000 13.805000 ;
        RECT 8.115000 13.805000 8.445000 13.845000 ;
        RECT 8.115000 13.845000 8.485000 13.885000 ;
        RECT 8.115000 13.885000 8.525000 13.975000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.785000 1.165000 65.565000 1.485000 ;
        RECT 65.110000 1.040000 65.565000 1.165000 ;
        RECT 65.235000 0.000000 65.565000 0.915000 ;
        RECT 65.235000 0.915000 65.565000 1.040000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.655000 0.000000 51.985000 7.760000 ;
        RECT 51.655000 7.760000 51.985000 7.910000 ;
        RECT 51.655000 7.910000 52.135000 8.060000 ;
        RECT 51.655000 8.060000 52.435000 8.380000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.105000 20.955000 129.435000 21.685000 ;
        RECT 129.125000  0.000000 129.455000 20.955000 ;
    END
  END DM[0]
  PIN DM[1]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.275000  0.000000 128.605000 19.875000 ;
        RECT 128.275000 19.875000 128.605000 19.885000 ;
        RECT 128.275000 19.885000 128.615000 19.895000 ;
        RECT 128.275000 19.895000 128.625000 20.180000 ;
        RECT 128.285000 20.180000 128.625000 20.190000 ;
        RECT 128.295000 20.190000 128.625000 20.200000 ;
        RECT 128.295000 20.200000 128.625000 21.685000 ;
    END
  END DM[1]
  PIN DM[2]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.375000 20.280000 108.725000 20.640000 ;
        RECT 108.375000 20.640000 108.705000 21.685000 ;
        RECT 108.395000  0.000000 108.725000 20.280000 ;
    END
  END DM[2]
  PIN ENABLE_H
    ANTENNAGATEAREA  8.880000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.135000  0.000000 22.465000 31.675000 ;
        RECT 22.135000 31.675000 22.465000 31.810000 ;
        RECT 22.135000 31.810000 22.600000 31.945000 ;
        RECT 22.135000 31.945000 22.875000 32.275000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.110000 0.000000 7.440000 19.735000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  3.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.770000 0.000000 9.100000 8.620000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    ANTENNAGATEAREA  6.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.845000 0.000000 96.215000 1.740000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    ANTENNAGATEAREA  3.120000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.765000 0.000000 6.365000 13.205000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    ANTENNAGATEAREA  1.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 19.635000  0.000000 19.965000 17.750000 ;
        RECT 19.635000 17.750000 19.965000 17.865000 ;
        RECT 19.635000 17.865000 20.080000 17.980000 ;
        RECT 19.635000 17.980000 20.195000 17.985000 ;
        RECT 19.675000 17.985000 20.200000 18.025000 ;
        RECT 19.715000 18.025000 20.240000 18.065000 ;
        RECT 19.830000 18.065000 20.280000 18.180000 ;
        RECT 19.945000 18.180000 20.280000 18.295000 ;
        RECT 19.950000 18.295000 20.280000 18.300000 ;
        RECT 19.950000 18.300000 20.280000 22.865000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.900000 14.055000 27.680000 14.375000 ;
        RECT 26.905000 14.050000 27.685000 14.055000 ;
        RECT 27.055000 13.900000 27.685000 14.050000 ;
        RECT 27.205000 13.750000 27.685000 13.900000 ;
        RECT 27.355000  0.000000 27.685000 13.600000 ;
        RECT 27.355000 13.600000 27.685000 13.750000 ;
    END
  END HLD_OVR
  PIN HYS_TRIM
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.905000 8.060000 45.685000 8.380000 ;
        RECT 45.055000 7.910000 45.685000 8.060000 ;
        RECT 45.205000 7.760000 45.685000 7.910000 ;
        RECT 45.355000 0.000000 45.685000 7.610000 ;
        RECT 45.355000 7.610000 45.685000 7.760000 ;
    END
  END HYS_TRIM
  PIN IB_MODE_SEL[0]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.815000 0.000000 87.145000 21.685000 ;
    END
  END IB_MODE_SEL[0]
  PIN IB_MODE_SEL[1]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.935000 0.000000 67.265000 21.685000 ;
    END
  END IB_MODE_SEL[1]
  PIN IN
    ANTENNAPARTIALMETALSIDEAREA  23.36800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.380000 0.000000 20.710000 15.275000 ;
    END
  END IN
  PIN INP_DIS
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.095000 8.060000 107.875000 8.380000 ;
        RECT 107.285000 8.055000 107.875000 8.060000 ;
        RECT 107.415000 7.925000 107.875000 8.055000 ;
        RECT 107.545000 0.000000 107.875000 7.795000 ;
        RECT 107.545000 7.795000 107.875000 7.925000 ;
    END
  END INP_DIS
  PIN IN_H
    ANTENNAPARTIALMETALSIDEAREA  1.722440 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.490000 0.610000 24.710000 0.940000 ;
        RECT 24.100000 0.605000 24.710000 0.610000 ;
        RECT 24.240000 0.465000 24.710000 0.605000 ;
        RECT 24.380000 0.000000 24.710000 0.325000 ;
        RECT 24.380000 0.325000 24.710000 0.465000 ;
    END
  END IN_H
  PIN OE_N
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.995000 8.060000 124.775000 8.380000 ;
        RECT 124.325000 7.940000 124.775000 8.060000 ;
        RECT 124.445000 0.000000 124.775000 7.820000 ;
        RECT 124.445000 7.820000 124.775000 7.940000 ;
    END
  END OE_N
  PIN OUT
    ANTENNAGATEAREA  1.529000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.125000  0.000000 74.455000 14.140000 ;
        RECT 74.125000 14.140000 74.455000 14.290000 ;
        RECT 74.125000 14.290000 74.605000 14.440000 ;
        RECT 74.125000 14.440000 74.755000 14.535000 ;
        RECT 74.125000 14.535000 78.505000 14.865000 ;
        RECT 77.870000 51.155000 78.600000 51.485000 ;
        RECT 77.930000 14.865000 78.505000 15.015000 ;
        RECT 77.950000 31.465000 78.355000 31.535000 ;
        RECT 77.950000 31.535000 78.285000 31.605000 ;
        RECT 77.950000 31.605000 78.280000 31.610000 ;
        RECT 77.950000 31.610000 78.280000 33.835000 ;
        RECT 77.950000 33.835000 78.280000 33.905000 ;
        RECT 77.950000 33.905000 78.350000 33.975000 ;
        RECT 77.950000 33.975000 78.420000 33.980000 ;
        RECT 77.990000 31.425000 78.425000 31.465000 ;
        RECT 77.990000 33.980000 78.425000 34.020000 ;
        RECT 78.030000 31.385000 78.465000 31.425000 ;
        RECT 78.030000 34.020000 78.465000 34.060000 ;
        RECT 78.035000 31.380000 78.505000 31.385000 ;
        RECT 78.080000 15.015000 78.505000 15.165000 ;
        RECT 78.100000 34.060000 78.505000 34.130000 ;
        RECT 78.105000 31.310000 78.505000 31.380000 ;
        RECT 78.170000 34.130000 78.505000 34.200000 ;
        RECT 78.175000 15.165000 78.505000 15.260000 ;
        RECT 78.175000 15.260000 78.505000 31.240000 ;
        RECT 78.175000 31.240000 78.505000 31.310000 ;
        RECT 78.175000 34.200000 78.505000 34.205000 ;
        RECT 78.175000 34.205000 78.505000 51.155000 ;
    END
  END OUT
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  228.2030 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 40.095000 132.705000 63.135000 147.730000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    ANTENNAPARTIALMETALSIDEAREA  256.0560 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.240000  5.465000 2.200000   5.470000 ;
        RECT 1.240000  5.470000 2.050000   5.620000 ;
        RECT 1.240000  5.620000 1.900000   5.770000 ;
        RECT 1.240000  5.770000 1.840000   5.830000 ;
        RECT 1.240000  5.830000 1.840000  70.535000 ;
        RECT 1.240000 70.535000 1.840000  70.680000 ;
        RECT 1.240000 70.680000 1.985000  70.825000 ;
        RECT 1.300000  5.405000 2.200000   5.465000 ;
        RECT 1.390000 70.825000 2.130000  70.975000 ;
        RECT 1.450000  5.255000 2.200000   5.405000 ;
        RECT 1.540000 70.975000 2.280000  71.125000 ;
        RECT 1.600000  0.000000 2.200000   5.105000 ;
        RECT 1.600000  5.105000 2.200000   5.255000 ;
        RECT 1.690000 71.125000 2.430000  71.275000 ;
        RECT 1.840000 71.275000 2.580000  71.425000 ;
        RECT 1.990000 71.425000 2.730000  71.575000 ;
        RECT 2.140000 71.575000 2.880000  71.725000 ;
        RECT 2.290000 71.725000 3.030000  71.875000 ;
        RECT 2.440000 71.875000 3.180000  72.025000 ;
        RECT 2.590000 72.025000 3.330000  72.175000 ;
        RECT 2.740000 72.175000 3.480000  72.325000 ;
        RECT 2.890000 72.325000 3.630000  72.475000 ;
        RECT 3.040000 72.475000 3.780000  72.625000 ;
        RECT 3.190000 72.625000 3.930000  72.775000 ;
        RECT 3.340000 72.775000 4.080000  72.925000 ;
        RECT 3.490000 72.925000 4.230000  73.075000 ;
        RECT 3.640000 73.075000 4.380000  73.225000 ;
        RECT 3.725000 73.225000 4.530000  73.310000 ;
        RECT 3.865000 73.310000 4.615000  73.450000 ;
        RECT 4.005000 73.450000 4.615000  73.590000 ;
        RECT 4.010000 73.590000 4.615000  73.595000 ;
        RECT 4.010000 73.595000 4.615000 159.560000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    ANTENNAPARTIALMETALSIDEAREA  257.9440 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.330000  0.000000 0.930000  71.100000 ;
        RECT 0.330000 71.100000 0.930000  71.240000 ;
        RECT 0.330000 71.240000 1.070000  71.380000 ;
        RECT 0.480000 71.380000 1.210000  71.530000 ;
        RECT 0.630000 71.530000 1.360000  71.680000 ;
        RECT 0.780000 71.680000 1.510000  71.830000 ;
        RECT 0.930000 71.830000 1.660000  71.980000 ;
        RECT 1.080000 71.980000 1.810000  72.130000 ;
        RECT 1.230000 72.130000 1.960000  72.280000 ;
        RECT 1.380000 72.280000 2.110000  72.430000 ;
        RECT 1.530000 72.430000 2.260000  72.580000 ;
        RECT 1.680000 72.580000 2.410000  72.730000 ;
        RECT 1.830000 72.730000 2.560000  72.880000 ;
        RECT 1.980000 72.880000 2.710000  73.030000 ;
        RECT 2.130000 73.030000 2.860000  73.180000 ;
        RECT 2.280000 73.180000 3.010000  73.330000 ;
        RECT 2.430000 73.330000 3.160000  73.480000 ;
        RECT 2.580000 73.480000 3.310000  73.630000 ;
        RECT 2.705000 73.630000 3.460000  73.755000 ;
        RECT 2.845000 73.755000 3.585000  73.895000 ;
        RECT 2.985000 73.895000 3.585000  74.035000 ;
        RECT 2.985000 74.035000 3.585000 160.945000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    ANTENNAPARTIALCUTAREA  0.120000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2.150000  6.260000 2.975000   6.410000 ;
        RECT 2.150000  6.410000 2.825000   6.560000 ;
        RECT 2.150000  6.560000 2.750000   6.635000 ;
        RECT 2.150000  6.635000 2.750000  70.075000 ;
        RECT 2.150000 70.075000 2.750000  70.220000 ;
        RECT 2.150000 70.220000 2.895000  70.365000 ;
        RECT 2.210000  6.200000 3.125000   6.260000 ;
        RECT 2.300000 70.365000 3.040000  70.515000 ;
        RECT 2.360000  6.050000 3.185000   6.200000 ;
        RECT 2.450000 70.515000 3.190000  70.665000 ;
        RECT 2.510000  5.900000 3.335000   6.050000 ;
        RECT 2.585000  5.825000 3.485000   5.900000 ;
        RECT 2.600000 70.665000 3.340000  70.815000 ;
        RECT 2.735000  5.675000 3.485000   5.825000 ;
        RECT 2.750000 70.815000 3.490000  70.965000 ;
        RECT 2.885000  0.000000 3.485000   5.525000 ;
        RECT 2.885000  5.525000 3.485000   5.675000 ;
        RECT 2.900000 70.965000 3.640000  71.115000 ;
        RECT 3.050000 71.115000 3.790000  71.265000 ;
        RECT 3.200000 71.265000 3.940000  71.415000 ;
        RECT 3.350000 71.415000 4.090000  71.565000 ;
        RECT 3.500000 71.565000 4.240000  71.715000 ;
        RECT 3.650000 71.715000 4.390000  71.865000 ;
        RECT 3.800000 71.865000 4.540000  72.015000 ;
        RECT 3.950000 72.015000 4.690000  72.165000 ;
        RECT 4.100000 72.165000 4.840000  72.315000 ;
        RECT 4.250000 72.315000 4.990000  72.465000 ;
        RECT 4.400000 72.465000 5.140000  72.615000 ;
        RECT 4.550000 72.615000 5.290000  72.765000 ;
        RECT 4.675000 72.765000 5.440000  72.890000 ;
        RECT 4.820000 72.890000 5.565000  73.035000 ;
        RECT 4.965000 73.035000 5.565000  73.180000 ;
        RECT 4.965000 73.180000 5.565000 122.920000 ;
    END
  END PAD_A_NOESD_H
  PIN SLEW_CTL[0]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.085000 0.000000 66.415000 21.685000 ;
    END
  END SLEW_CTL[0]
  PIN SLEW_CTL[1]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.205000 0.000000 46.535000 21.685000 ;
    END
  END SLEW_CTL[1]
  PIN SLOW
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 124.580000 12.150000 125.135000 12.300000 ;
        RECT 124.580000 12.300000 124.985000 12.450000 ;
        RECT 124.580000 12.450000 124.910000 12.525000 ;
        RECT 124.580000 12.525000 124.910000 18.470000 ;
        RECT 124.580000 18.470000 124.910000 18.615000 ;
        RECT 124.580000 18.615000 125.055000 18.760000 ;
        RECT 124.580000 18.760000 125.200000 18.765000 ;
        RECT 124.585000 12.145000 125.285000 12.150000 ;
        RECT 124.675000 12.055000 125.290000 12.145000 ;
        RECT 124.710000 18.765000 125.205000 18.895000 ;
        RECT 124.765000 11.965000 125.380000 12.055000 ;
        RECT 124.840000 11.890000 125.470000 11.965000 ;
        RECT 124.840000 18.895000 125.335000 19.025000 ;
        RECT 124.845000 19.025000 125.465000 19.030000 ;
        RECT 124.990000 11.740000 125.470000 11.890000 ;
        RECT 124.990000 19.030000 125.470000 19.175000 ;
        RECT 125.135000 19.175000 125.470000 19.320000 ;
        RECT 125.140000  0.000000 125.470000 11.590000 ;
        RECT 125.140000 11.590000 125.470000 11.740000 ;
        RECT 125.140000 19.320000 125.470000 19.325000 ;
        RECT 125.140000 19.325000 125.470000 31.390000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    ANTENNAGATEAREA 21 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.975000   0.000000 130.305000  61.465000 ;
        RECT 129.975000  61.465000 130.305000  61.560000 ;
        RECT 129.975000  61.560000 130.400000  61.655000 ;
        RECT 130.125000  61.655000 130.495000  61.805000 ;
        RECT 130.275000  61.805000 130.645000  61.955000 ;
        RECT 130.425000  61.955000 130.795000  62.105000 ;
        RECT 130.460000 110.205000 131.140000 110.935000 ;
        RECT 130.575000  62.105000 130.945000  62.255000 ;
        RECT 130.620000  62.255000 131.095000  62.300000 ;
        RECT 130.715000  62.300000 131.140000  62.395000 ;
        RECT 130.730000 110.125000 131.140000 110.205000 ;
        RECT 130.810000  62.395000 131.140000  62.490000 ;
        RECT 130.810000  62.490000 131.140000 110.045000 ;
        RECT 130.810000 110.045000 131.140000 110.125000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 114.650000 111.180000 115.485000 111.265000 ;
        RECT 114.650000 111.265000 115.400000 111.350000 ;
        RECT 114.670000 111.160000 115.570000 111.180000 ;
        RECT 114.820000 111.010000 115.590000 111.160000 ;
        RECT 114.970000 110.860000 115.740000 111.010000 ;
        RECT 114.990000 110.840000 115.890000 110.860000 ;
        RECT 115.140000 110.690000 115.890000 110.840000 ;
        RECT 115.290000   0.000000 115.890000 110.540000 ;
        RECT 115.290000 110.540000 115.890000 110.690000 ;
    END
  END TIE_LO_ESD
  PIN VINREF
    ANTENNAGATEAREA 54 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.035000 0.000000 44.365000 4.460000 ;
        RECT 44.035000 4.460000 44.365000 4.610000 ;
        RECT 44.035000 4.610000 44.515000 4.760000 ;
        RECT 44.035000 4.760000 44.665000 4.860000 ;
        RECT 44.035000 4.860000 44.765000 5.190000 ;
    END
  END VINREF
  PIN VTRIP_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.665000 0.000000 87.995000 21.685000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.255000  8.930000 140.000000 13.465000 ;
        RECT 138.730000  8.885000 140.000000  8.930000 ;
        RECT 138.730000 13.465000 140.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 8.985000 140.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 2.035000 140.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 2.135000 140.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.035000 14.935000 140.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 139.035000 15.035000 140.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 19.785000 140.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 70.035000 140.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 19.885000 140.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 70.035000 140.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 64.085000 140.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 64.185000 140.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 36.735000 140.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 47.735000 140.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 51.645000 140.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 56.405000 140.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 36.840000 140.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 47.735000 140.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 41.585000 140.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 41.685000 140.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 175.785000 140.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 25.835000 140.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 175.785000 140.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 25.935000 140.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 58.235000 140.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 58.335000 140.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730000 31.885000 140.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730000 31.985000 140.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  10.485000 187.010000  10.715000 187.105000 ;
      RECT  10.485000 187.105000  10.830000 187.335000 ;
      RECT  11.220000 170.660000  15.760000 172.700000 ;
      RECT  11.395000 162.715000  13.005000 163.245000 ;
      RECT  11.600000  17.150000  16.580000  18.770000 ;
      RECT  11.600000  18.770000 140.000000  20.300000 ;
      RECT  11.600000  20.300000  22.570000  20.755000 ;
      RECT  13.915000 162.715000  15.525000 163.245000 ;
      RECT  18.005000  10.045000  18.175000  10.575000 ;
      RECT  32.245000  17.150000 140.000000  18.770000 ;
      RECT  69.500000  59.375000  69.820000  59.965000 ;
      RECT  84.135000  47.800000  88.065000  47.970000 ;
      RECT 118.305000 114.495000 140.145000 116.765000 ;
      RECT 120.645000  82.020000 123.195000  96.125000 ;
      RECT 120.725000  81.690000 123.195000  82.020000 ;
      RECT 129.625000  57.445000 131.645000  58.925000 ;
      RECT 131.375000 110.400000 140.145000 114.495000 ;
      RECT 135.060000  74.915000 135.565000 104.150000 ;
      RECT 135.140000  74.890000 135.565000  74.915000 ;
      RECT 135.140000 104.150000 135.565000 104.230000 ;
      RECT 136.065000 186.065000 138.125000 186.295000 ;
      RECT 136.065000 186.295000 136.295000 186.895000 ;
      RECT 136.065000 187.570000 136.295000 187.870000 ;
      RECT 136.065000 187.870000 138.125000 188.100000 ;
      RECT 136.815000 187.175000 137.345000 187.345000 ;
      RECT 137.895000 186.295000 138.125000 187.870000 ;
    LAYER met1 ;
      RECT   0.000000  0.000000 140.000000 200.000000 ;
      RECT 140.000000 53.225000 140.350000  53.955000 ;
      RECT 140.000000 63.715000 140.160000  64.685000 ;
    LAYER met2 ;
      RECT 0.000000  0.000000 140.000000  63.715000 ;
      RECT 0.000000 63.715000 140.325000  68.140000 ;
      RECT 0.000000 68.140000 140.000000 200.000000 ;
    LAYER met3 ;
      RECT   0.000000   0.000000   0.030000  71.505000 ;
      RECT   0.000000  71.505000   2.685000  74.160000 ;
      RECT   0.000000  71.765000   0.150000  71.915000 ;
      RECT   0.000000  71.915000   0.300000  72.065000 ;
      RECT   0.000000  72.065000   0.450000  72.215000 ;
      RECT   0.000000  72.215000   0.600000  72.365000 ;
      RECT   0.000000  72.365000   0.750000  72.515000 ;
      RECT   0.000000  72.515000   0.900000  72.665000 ;
      RECT   0.000000  72.665000   1.050000  72.815000 ;
      RECT   0.000000  72.815000   1.200000  72.965000 ;
      RECT   0.000000  72.965000   1.350000  73.115000 ;
      RECT   0.000000  73.115000   1.500000  73.265000 ;
      RECT   0.000000  73.265000   1.650000  73.415000 ;
      RECT   0.000000  73.415000   1.800000  73.565000 ;
      RECT   0.000000  73.565000   1.950000  73.715000 ;
      RECT   0.000000  73.715000   2.100000  73.865000 ;
      RECT   0.000000  73.865000   2.250000  74.015000 ;
      RECT   0.000000  74.015000   2.400000  74.165000 ;
      RECT   0.000000  74.160000   2.685000 161.245000 ;
      RECT   0.000000  74.165000   2.550000  74.200000 ;
      RECT   0.000000  74.200000   2.585000 161.345000 ;
      RECT   0.000000 161.245000 140.000000 200.000000 ;
      RECT   0.000000 161.345000 140.000000 200.000000 ;
      RECT   1.230000   0.000000   1.300000   4.980000 ;
      RECT   2.500000   0.000000   2.585000   5.400000 ;
      RECT   3.050000   6.760000   5.465000  13.505000 ;
      RECT   3.050000  13.505000   6.810000  20.035000 ;
      RECT   3.050000  20.035000  19.650000  23.165000 ;
      RECT   3.050000  23.165000  21.835000  32.575000 ;
      RECT   3.050000  32.575000  77.650000  34.105000 ;
      RECT   3.050000  34.105000  77.875000  34.330000 ;
      RECT   3.050000  34.330000  77.875000  50.855000 ;
      RECT   3.050000  50.855000  77.570000  51.785000 ;
      RECT   3.050000  51.785000 114.990000  69.950000 ;
      RECT   3.050000  69.950000 114.990000  72.765000 ;
      RECT   3.150000   6.800000   5.365000  13.605000 ;
      RECT   3.150000  13.605000   6.710000  20.135000 ;
      RECT   3.150000  13.605000   6.710000  23.265000 ;
      RECT   3.150000  20.135000  19.550000  23.265000 ;
      RECT   3.150000  20.135000  19.550000  32.675000 ;
      RECT   3.150000  23.265000  21.735000  32.675000 ;
      RECT   3.150000  23.265000  21.735000  34.145000 ;
      RECT   3.150000  23.265000  21.735000  34.145000 ;
      RECT   3.150000  23.265000  21.735000  34.145000 ;
      RECT   3.150000  32.675000  77.550000  34.145000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  32.675000  77.550000  50.755000 ;
      RECT   3.150000  34.145000  77.550000  34.260000 ;
      RECT   3.150000  34.145000  77.550000  34.260000 ;
      RECT   3.150000  34.260000  77.665000  34.370000 ;
      RECT   3.150000  34.260000  77.665000  34.370000 ;
      RECT   3.150000  34.370000  77.470000  51.885000 ;
      RECT   3.150000  34.370000  77.470000  69.910000 ;
      RECT   3.150000  34.370000  77.775000  50.755000 ;
      RECT   3.150000  50.755000  77.470000  51.885000 ;
      RECT   3.150000  51.885000 114.890000  69.910000 ;
      RECT   3.285000   6.665000   5.365000   6.800000 ;
      RECT   3.300000  69.910000 114.890000  70.060000 ;
      RECT   3.300000  69.910000 114.890000  70.060000 ;
      RECT   3.435000   6.515000   5.365000   6.665000 ;
      RECT   3.450000  70.060000 114.890000  70.210000 ;
      RECT   3.450000  70.060000 114.890000  70.210000 ;
      RECT   3.585000   6.365000   5.365000   6.515000 ;
      RECT   3.600000  70.210000 114.890000  70.360000 ;
      RECT   3.600000  70.210000 114.890000  70.360000 ;
      RECT   3.735000   6.215000   5.365000   6.365000 ;
      RECT   3.750000  70.360000 114.890000  70.510000 ;
      RECT   3.750000  70.360000 114.890000  70.510000 ;
      RECT   3.785000   0.000000   5.465000   6.025000 ;
      RECT   3.785000   6.025000   5.465000   6.760000 ;
      RECT   3.885000   0.000000   5.365000   6.065000 ;
      RECT   3.885000   6.065000   5.365000   6.215000 ;
      RECT   3.885000 159.860000 140.000000 161.245000 ;
      RECT   3.900000  70.510000 114.890000  70.660000 ;
      RECT   3.900000  70.510000 114.890000  70.660000 ;
      RECT   3.985000 159.960000 140.000000 161.345000 ;
      RECT   3.985000 159.960000 140.000000 200.000000 ;
      RECT   4.050000  70.660000 114.890000  70.810000 ;
      RECT   4.050000  70.660000 114.890000  70.810000 ;
      RECT   4.200000  70.810000 114.890000  70.960000 ;
      RECT   4.200000  70.810000 114.890000  70.960000 ;
      RECT   4.350000  70.960000 114.890000  71.110000 ;
      RECT   4.350000  70.960000 114.890000  71.110000 ;
      RECT   4.500000  71.110000 114.890000  71.260000 ;
      RECT   4.500000  71.110000 114.890000  71.260000 ;
      RECT   4.650000  71.260000 114.890000  71.410000 ;
      RECT   4.650000  71.260000 114.890000  71.410000 ;
      RECT   4.800000  71.410000 114.890000  71.560000 ;
      RECT   4.800000  71.410000 114.890000  71.560000 ;
      RECT   4.915000 123.220000 140.000000 159.860000 ;
      RECT   4.950000  71.560000 114.890000  71.710000 ;
      RECT   4.950000  71.560000 114.890000  71.710000 ;
      RECT   5.015000 123.320000 140.000000 159.960000 ;
      RECT   5.015000 123.320000 140.000000 200.000000 ;
      RECT   5.100000  71.710000 114.890000  71.860000 ;
      RECT   5.100000  71.710000 114.890000  71.860000 ;
      RECT   5.250000  71.860000 114.890000  72.010000 ;
      RECT   5.250000  71.860000 114.890000  72.010000 ;
      RECT   5.400000  72.010000 114.890000  72.160000 ;
      RECT   5.400000  72.010000 114.890000  72.160000 ;
      RECT   5.550000  72.160000 114.890000  72.310000 ;
      RECT   5.550000  72.160000 114.890000  72.310000 ;
      RECT   5.700000  72.310000 114.890000  72.460000 ;
      RECT   5.700000  72.310000 114.890000  72.460000 ;
      RECT   5.850000  72.460000 114.890000  72.610000 ;
      RECT   5.850000  72.460000 114.890000  72.610000 ;
      RECT   5.865000  72.765000 114.990000 110.415000 ;
      RECT   5.865000 110.415000 114.350000 111.055000 ;
      RECT   5.865000 111.055000 114.350000 111.650000 ;
      RECT   5.865000 111.650000 114.965000 112.210000 ;
      RECT   5.865000 112.210000 140.000000 123.220000 ;
      RECT   5.965000  72.610000 114.890000  72.725000 ;
      RECT   5.965000  72.610000 114.890000  72.725000 ;
      RECT   5.965000  72.725000 114.890000 110.375000 ;
      RECT   5.965000 110.375000 114.250000 123.320000 ;
      RECT   5.965000 110.375000 114.250000 123.320000 ;
      RECT   5.965000 110.375000 114.250000 123.320000 ;
      RECT   5.965000 110.375000 114.740000 110.525000 ;
      RECT   5.965000 110.375000 114.740000 110.525000 ;
      RECT   5.965000 110.525000 114.590000 110.675000 ;
      RECT   5.965000 110.525000 114.590000 110.675000 ;
      RECT   5.965000 110.675000 114.440000 110.825000 ;
      RECT   5.965000 110.675000 114.440000 110.825000 ;
      RECT   5.965000 110.825000 114.290000 110.975000 ;
      RECT   5.965000 110.825000 114.290000 110.975000 ;
      RECT   5.965000 110.975000 114.250000 111.015000 ;
      RECT   5.965000 110.975000 114.250000 111.015000 ;
      RECT   5.965000 111.015000 114.250000 111.750000 ;
      RECT   5.965000 111.750000 114.865000 112.450000 ;
      RECT   5.965000 111.750000 114.865000 123.320000 ;
      RECT   5.965000 111.750000 114.865000 123.320000 ;
      RECT   5.965000 111.750000 114.865000 123.320000 ;
      RECT   5.965000 112.450000 140.000000 123.320000 ;
      RECT   6.665000   0.000000   6.810000  13.505000 ;
      RECT   7.740000   0.000000   7.815000  13.760000 ;
      RECT   7.740000  14.690000  19.335000  18.110000 ;
      RECT   7.740000  18.110000  19.650000  18.425000 ;
      RECT   7.740000  18.425000  19.650000  20.035000 ;
      RECT   7.840000  14.790000  19.235000  18.150000 ;
      RECT   7.840000  14.790000  19.235000  18.465000 ;
      RECT   7.840000  18.150000  19.235000  18.300000 ;
      RECT   7.840000  18.150000  19.235000  18.300000 ;
      RECT   7.840000  18.300000  19.385000  18.450000 ;
      RECT   7.840000  18.300000  19.385000  18.450000 ;
      RECT   7.840000  18.450000  19.535000  18.465000 ;
      RECT   7.840000  18.450000  19.535000  18.465000 ;
      RECT   7.840000  18.465000  19.550000  20.135000 ;
      RECT   7.840000  18.465000  19.550000  32.675000 ;
      RECT   8.745000   8.920000  19.335000  13.680000 ;
      RECT   8.745000  13.680000  19.335000  13.945000 ;
      RECT   8.845000   9.020000  19.235000  13.640000 ;
      RECT   8.975000  13.640000  19.235000  13.770000 ;
      RECT   8.975000  13.640000  19.235000  13.770000 ;
      RECT   9.010000  13.945000  19.335000  14.690000 ;
      RECT   9.105000  13.770000  19.235000  13.900000 ;
      RECT   9.105000  13.770000  19.235000  13.900000 ;
      RECT   9.110000   9.020000  19.235000  18.150000 ;
      RECT   9.110000  13.900000  19.235000  13.905000 ;
      RECT   9.110000  13.900000  19.235000  13.905000 ;
      RECT   9.110000  13.905000  19.235000  14.790000 ;
      RECT   9.400000   0.000000  19.335000   8.920000 ;
      RECT   9.500000   0.000000  19.235000   9.020000 ;
      RECT  20.265000  15.575000  21.835000  17.625000 ;
      RECT  20.265000  17.625000  21.835000  17.940000 ;
      RECT  20.365000  15.675000  21.735000  17.585000 ;
      RECT  20.515000  17.585000  21.735000  17.735000 ;
      RECT  20.580000  17.940000  21.835000  23.165000 ;
      RECT  20.665000  17.735000  21.735000  17.885000 ;
      RECT  20.680000  17.885000  21.735000  17.900000 ;
      RECT  20.680000  17.900000  21.735000  23.265000 ;
      RECT  21.010000   0.000000  21.835000  15.575000 ;
      RECT  21.110000   0.000000  21.735000  15.675000 ;
      RECT  22.765000   0.000000  24.080000   0.200000 ;
      RECT  22.765000   0.200000  23.970000   0.310000 ;
      RECT  22.765000   0.310000  23.190000   1.240000 ;
      RECT  22.765000   1.240000  27.055000  13.475000 ;
      RECT  22.765000  13.475000  26.600000  13.930000 ;
      RECT  22.765000  13.930000  26.600000  14.675000 ;
      RECT  22.765000  14.675000  45.905000  21.985000 ;
      RECT  22.765000  21.985000  77.875000  31.115000 ;
      RECT  22.765000  31.115000  77.650000  31.340000 ;
      RECT  22.765000  31.340000  77.650000  31.550000 ;
      RECT  22.765000  31.550000  77.650000  31.645000 ;
      RECT  22.865000   1.340000  26.955000  13.435000 ;
      RECT  22.865000  13.435000  26.500000  22.085000 ;
      RECT  22.865000  13.435000  26.500000  22.085000 ;
      RECT  22.865000  13.435000  26.805000  13.585000 ;
      RECT  22.865000  13.435000  26.805000  13.585000 ;
      RECT  22.865000  13.585000  26.655000  13.735000 ;
      RECT  22.865000  13.585000  26.655000  13.735000 ;
      RECT  22.865000  13.735000  26.505000  13.885000 ;
      RECT  22.865000  13.735000  26.505000  13.885000 ;
      RECT  22.865000  13.885000  26.500000  13.890000 ;
      RECT  22.865000  13.885000  26.500000  13.890000 ;
      RECT  22.865000  13.890000  26.500000  14.775000 ;
      RECT  22.865000  14.775000  45.805000  22.085000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.550000  31.545000 ;
      RECT  22.865000  22.085000  77.775000  31.075000 ;
      RECT  22.865000  31.075000  77.665000  31.185000 ;
      RECT  22.865000  31.075000  77.665000  31.185000 ;
      RECT  22.865000  31.185000  77.555000  31.295000 ;
      RECT  22.865000  31.185000  77.555000  31.295000 ;
      RECT  22.865000  31.295000  77.550000  31.300000 ;
      RECT  22.865000  31.295000  77.550000  31.300000 ;
      RECT  22.865000  31.300000  77.550000  31.545000 ;
      RECT  23.175000  31.645000  77.650000  32.575000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  22.085000  77.550000  50.755000 ;
      RECT  23.275000  31.545000  77.550000  32.675000 ;
      RECT  25.010000   0.000000  27.055000   1.240000 ;
      RECT  25.110000   0.000000  26.955000   1.340000 ;
      RECT  27.980000  14.355000  45.905000  14.675000 ;
      RECT  27.985000   0.000000  43.735000   5.490000 ;
      RECT  27.985000   5.490000  45.055000   7.485000 ;
      RECT  27.985000   7.485000  44.605000   7.935000 ;
      RECT  27.985000   7.935000  44.605000   8.680000 ;
      RECT  27.985000   8.680000  45.905000  14.355000 ;
      RECT  28.080000  14.455000  45.805000  14.775000 ;
      RECT  28.080000  14.455000  45.805000  22.085000 ;
      RECT  28.085000   0.000000  43.635000   5.590000 ;
      RECT  28.085000   0.000000  43.635000  14.455000 ;
      RECT  28.085000   0.000000  43.635000  14.455000 ;
      RECT  28.085000   5.590000  44.505000  14.455000 ;
      RECT  28.085000   5.590000  44.505000  14.455000 ;
      RECT  28.085000   5.590000  44.955000   7.445000 ;
      RECT  28.085000   7.445000  44.805000   7.595000 ;
      RECT  28.085000   7.445000  44.805000   7.595000 ;
      RECT  28.085000   7.595000  44.655000   7.745000 ;
      RECT  28.085000   7.595000  44.655000   7.745000 ;
      RECT  28.085000   7.745000  44.505000   7.895000 ;
      RECT  28.085000   7.745000  44.505000   7.895000 ;
      RECT  28.085000   7.895000  44.505000   8.780000 ;
      RECT  28.085000   8.780000  45.805000  14.455000 ;
      RECT  28.085000   8.780000  45.805000  14.775000 ;
      RECT  28.085000   8.780000  45.805000  22.085000 ;
      RECT  44.665000   0.000000  45.055000   4.335000 ;
      RECT  44.665000   4.335000  45.055000   4.725000 ;
      RECT  46.835000   0.000000  51.355000   8.680000 ;
      RECT  46.835000   8.680000  65.785000  21.985000 ;
      RECT  46.935000   0.000000  51.255000   8.780000 ;
      RECT  46.935000   0.000000  51.255000  22.085000 ;
      RECT  46.935000   0.000000  51.255000  22.085000 ;
      RECT  46.935000   0.000000  51.255000  22.085000 ;
      RECT  46.935000   8.780000  65.685000  22.085000 ;
      RECT  52.285000   0.000000  64.935000   0.790000 ;
      RECT  52.285000   0.790000  64.860000   0.865000 ;
      RECT  52.285000   0.865000  64.485000   1.785000 ;
      RECT  52.285000   1.785000  65.785000   7.635000 ;
      RECT  52.285000   7.635000  65.785000   7.760000 ;
      RECT  52.385000   0.000000  64.835000   0.765000 ;
      RECT  52.385000   0.765000  64.385000   3.005000 ;
      RECT  52.385000   1.885000  65.685000   7.660000 ;
      RECT  52.735000   7.760000  65.785000   8.680000 ;
      RECT  52.835000   1.885000  65.685000  22.085000 ;
      RECT  52.835000   7.660000  65.685000   8.780000 ;
      RECT  67.565000   0.000000  73.825000  15.165000 ;
      RECT  67.565000  15.165000  77.875000  15.385000 ;
      RECT  67.565000  15.385000  77.875000  21.985000 ;
      RECT  67.665000   0.000000  73.725000  15.265000 ;
      RECT  67.665000  15.265000  77.615000  15.345000 ;
      RECT  67.665000  15.265000  77.615000  15.345000 ;
      RECT  67.665000  15.345000  77.695000  15.425000 ;
      RECT  67.665000  15.345000  77.695000  15.425000 ;
      RECT  67.665000  15.425000  77.775000  22.085000 ;
      RECT  74.755000   0.000000  86.515000  14.015000 ;
      RECT  74.755000  14.015000  86.515000  14.235000 ;
      RECT  74.855000   0.000000  86.510000  13.975000 ;
      RECT  74.935000  13.975000  86.510000  14.055000 ;
      RECT  74.935000  13.975000  86.510000  14.055000 ;
      RECT  75.015000  14.055000  86.510000  14.135000 ;
      RECT  75.015000  14.055000  86.510000  14.135000 ;
      RECT  78.580000  31.735000 114.990000  33.710000 ;
      RECT  78.580000  33.710000 114.990000  33.935000 ;
      RECT  78.680000  31.775000 114.890000  33.670000 ;
      RECT  78.790000  31.665000 114.890000  31.775000 ;
      RECT  78.790000  31.665000 114.890000  31.775000 ;
      RECT  78.790000  33.670000 114.890000  33.780000 ;
      RECT  78.790000  33.670000 114.890000  33.780000 ;
      RECT  78.805000  14.235000  86.515000  21.985000 ;
      RECT  78.805000  21.985000 114.990000  31.510000 ;
      RECT  78.805000  31.510000 114.990000  31.735000 ;
      RECT  78.805000  33.935000 114.990000  50.855000 ;
      RECT  78.900000  33.780000 114.890000  33.890000 ;
      RECT  78.900000  33.780000 114.890000  33.890000 ;
      RECT  78.900000  50.855000 114.990000  51.785000 ;
      RECT  78.905000  14.135000  86.510000  22.085000 ;
      RECT  78.905000  14.135000  86.510000  31.550000 ;
      RECT  78.905000  22.085000 114.890000  31.550000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  22.085000 114.890000  33.895000 ;
      RECT  78.905000  31.550000 114.890000  31.665000 ;
      RECT  78.905000  31.550000 114.890000  31.665000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.670000 114.890000  50.755000 ;
      RECT  78.905000  33.890000 114.890000  33.895000 ;
      RECT  78.905000  33.890000 114.890000  33.895000 ;
      RECT  78.905000  33.895000 114.890000  50.755000 ;
      RECT  79.000000  33.895000 114.890000  69.910000 ;
      RECT  79.000000  33.895000 114.890000  69.910000 ;
      RECT  79.000000  50.755000 114.890000  51.885000 ;
      RECT  88.295000   0.000000  95.545000   2.040000 ;
      RECT  88.295000   2.040000 107.245000   7.670000 ;
      RECT  88.295000   7.670000 107.155000   7.760000 ;
      RECT  88.295000   7.760000 106.795000   8.680000 ;
      RECT  88.295000   8.680000 108.095000  19.980000 ;
      RECT  88.295000  19.980000 108.075000  21.985000 ;
      RECT  88.395000   0.000000  95.445000   2.140000 ;
      RECT  88.395000   0.000000  95.445000   7.660000 ;
      RECT  88.395000   0.000000  95.445000   7.660000 ;
      RECT  88.395000   2.140000 106.695000  19.880000 ;
      RECT  88.395000   2.140000 107.145000   7.660000 ;
      RECT  88.395000   7.660000 106.695000   8.780000 ;
      RECT  88.395000   8.780000 107.975000  22.085000 ;
      RECT  88.395000   8.780000 107.975000  22.085000 ;
      RECT  88.395000   8.780000 107.995000  19.880000 ;
      RECT  88.395000  19.880000 107.975000  22.085000 ;
      RECT  96.515000   0.000000 107.245000   2.040000 ;
      RECT  96.615000   0.000000 107.145000   2.140000 ;
      RECT  96.615000   0.000000 107.145000   7.660000 ;
      RECT  96.615000   0.000000 107.145000   7.660000 ;
      RECT 109.005000  20.940000 114.990000  21.985000 ;
      RECT 109.025000   0.000000 114.990000  20.940000 ;
      RECT 109.105000  21.040000 114.890000  22.085000 ;
      RECT 109.125000   0.000000 114.890000  21.040000 ;
      RECT 109.125000   0.000000 114.890000  22.085000 ;
      RECT 109.125000   0.000000 114.890000  22.085000 ;
      RECT 114.930000 112.385000 140.000000 112.450000 ;
      RECT 114.930000 112.385000 140.000000 112.450000 ;
      RECT 115.080000 112.235000 140.000000 112.385000 ;
      RECT 115.080000 112.235000 140.000000 112.385000 ;
      RECT 115.230000 112.085000 140.000000 112.235000 ;
      RECT 115.230000 112.085000 140.000000 112.235000 ;
      RECT 115.380000 111.935000 140.000000 112.085000 ;
      RECT 115.380000 111.935000 140.000000 112.085000 ;
      RECT 115.530000 111.785000 140.000000 111.935000 ;
      RECT 115.530000 111.785000 140.000000 111.935000 ;
      RECT 115.680000 111.635000 140.000000 111.785000 ;
      RECT 115.680000 111.635000 140.000000 111.785000 ;
      RECT 115.830000 111.485000 140.000000 111.635000 ;
      RECT 115.830000 111.485000 140.000000 111.635000 ;
      RECT 115.940000 111.235000 140.000000 112.210000 ;
      RECT 115.980000 111.335000 140.000000 111.485000 ;
      RECT 115.980000 111.335000 140.000000 111.485000 ;
      RECT 115.990000 111.325000 130.060000 111.335000 ;
      RECT 115.990000 111.325000 130.060000 111.335000 ;
      RECT 116.140000 111.175000 130.060000 111.325000 ;
      RECT 116.140000 111.175000 130.060000 111.325000 ;
      RECT 116.190000   0.000000 124.145000   7.695000 ;
      RECT 116.190000   7.695000 124.080000   7.760000 ;
      RECT 116.190000   7.760000 123.695000   8.680000 ;
      RECT 116.190000   8.680000 124.840000  11.465000 ;
      RECT 116.190000  11.465000 124.280000  12.025000 ;
      RECT 116.190000  12.025000 124.280000  18.890000 ;
      RECT 116.190000  18.890000 124.840000  19.450000 ;
      RECT 116.190000  19.450000 124.840000  31.690000 ;
      RECT 116.190000  31.690000 129.675000  61.780000 ;
      RECT 116.190000  61.780000 130.510000  62.615000 ;
      RECT 116.190000  62.615000 130.510000 109.905000 ;
      RECT 116.190000 109.905000 130.160000 110.985000 ;
      RECT 116.190000 110.985000 130.160000 111.235000 ;
      RECT 116.290000   0.000000 123.595000  11.985000 ;
      RECT 116.290000   0.000000 123.595000  18.930000 ;
      RECT 116.290000   0.000000 124.045000   7.660000 ;
      RECT 116.290000   7.660000 123.595000   8.780000 ;
      RECT 116.290000   8.780000 124.180000  18.930000 ;
      RECT 116.290000   8.780000 124.740000  11.425000 ;
      RECT 116.290000  11.425000 124.590000  11.575000 ;
      RECT 116.290000  11.425000 124.590000  11.575000 ;
      RECT 116.290000  11.575000 124.440000  11.725000 ;
      RECT 116.290000  11.575000 124.440000  11.725000 ;
      RECT 116.290000  11.725000 124.290000  11.875000 ;
      RECT 116.290000  11.725000 124.290000  11.875000 ;
      RECT 116.290000  11.875000 124.180000  11.985000 ;
      RECT 116.290000  11.875000 124.180000  11.985000 ;
      RECT 116.290000  11.985000 124.180000  18.930000 ;
      RECT 116.290000  11.985000 124.180000  19.490000 ;
      RECT 116.290000  18.930000 124.180000  19.080000 ;
      RECT 116.290000  18.930000 124.180000  19.080000 ;
      RECT 116.290000  19.080000 124.330000  19.230000 ;
      RECT 116.290000  19.080000 124.330000  19.230000 ;
      RECT 116.290000  19.230000 124.480000  19.380000 ;
      RECT 116.290000  19.230000 124.480000  19.380000 ;
      RECT 116.290000  19.380000 124.630000  19.490000 ;
      RECT 116.290000  19.380000 124.630000  19.490000 ;
      RECT 116.290000  19.490000 124.740000  31.790000 ;
      RECT 116.290000  19.490000 124.740000  61.820000 ;
      RECT 116.290000  31.790000 129.575000  61.820000 ;
      RECT 116.290000  61.820000 129.575000  61.970000 ;
      RECT 116.290000  61.820000 129.575000  61.970000 ;
      RECT 116.290000  61.970000 129.725000  62.120000 ;
      RECT 116.290000  61.970000 129.725000  62.120000 ;
      RECT 116.290000  62.120000 129.875000  62.270000 ;
      RECT 116.290000  62.120000 129.875000  62.270000 ;
      RECT 116.290000  62.270000 130.025000  62.420000 ;
      RECT 116.290000  62.270000 130.025000  62.420000 ;
      RECT 116.290000  62.420000 130.175000  62.570000 ;
      RECT 116.290000  62.420000 130.175000  62.570000 ;
      RECT 116.290000  62.570000 130.325000  62.655000 ;
      RECT 116.290000  62.570000 130.325000  62.655000 ;
      RECT 116.290000  62.655000 130.410000 109.805000 ;
      RECT 116.290000 109.805000 130.060000 111.025000 ;
      RECT 116.290000 111.025000 130.060000 111.175000 ;
      RECT 116.290000 111.025000 130.060000 111.175000 ;
      RECT 125.210000  12.650000 127.975000  18.345000 ;
      RECT 125.210000  18.345000 127.975000  18.905000 ;
      RECT 125.310000  12.690000 127.875000  18.305000 ;
      RECT 125.420000  12.580000 127.875000  12.690000 ;
      RECT 125.460000  18.305000 127.875000  18.455000 ;
      RECT 125.570000  12.430000 127.875000  12.580000 ;
      RECT 125.610000  18.455000 127.875000  18.605000 ;
      RECT 125.720000  12.280000 127.875000  12.430000 ;
      RECT 125.760000  18.605000 127.875000  18.755000 ;
      RECT 125.770000   0.000000 127.975000  12.090000 ;
      RECT 125.770000  12.090000 127.975000  12.650000 ;
      RECT 125.770000  18.905000 127.975000  20.305000 ;
      RECT 125.770000  20.305000 127.995000  20.325000 ;
      RECT 125.770000  20.325000 127.995000  21.985000 ;
      RECT 125.770000  21.985000 129.675000  31.690000 ;
      RECT 125.870000   0.000000 127.875000  12.130000 ;
      RECT 125.870000  12.130000 127.875000  12.280000 ;
      RECT 125.870000  18.755000 127.875000  18.865000 ;
      RECT 125.870000  18.865000 127.875000  20.345000 ;
      RECT 125.870000  20.345000 127.875000  20.355000 ;
      RECT 125.870000  20.355000 127.885000  20.365000 ;
      RECT 125.870000  20.365000 127.895000  22.085000 ;
      RECT 125.870000  22.085000 129.575000  31.790000 ;
      RECT 130.605000   0.000000 140.000000  61.340000 ;
      RECT 130.605000  61.340000 140.000000  62.175000 ;
      RECT 130.705000   0.000000 140.000000  61.300000 ;
      RECT 130.855000  61.300000 140.000000  61.450000 ;
      RECT 130.855000  61.300000 140.000000  61.450000 ;
      RECT 131.005000  61.450000 140.000000  61.600000 ;
      RECT 131.005000  61.450000 140.000000  61.600000 ;
      RECT 131.155000  61.600000 140.000000  61.750000 ;
      RECT 131.155000  61.600000 140.000000  61.750000 ;
      RECT 131.305000  61.750000 140.000000  61.900000 ;
      RECT 131.305000  61.750000 140.000000  61.900000 ;
      RECT 131.440000  62.175000 140.000000 111.235000 ;
      RECT 131.455000  61.900000 140.000000  62.050000 ;
      RECT 131.455000  61.900000 140.000000  62.050000 ;
      RECT 131.540000  62.050000 140.000000  62.135000 ;
      RECT 131.540000  62.050000 140.000000  62.135000 ;
      RECT 131.540000  62.135000 140.000000 111.335000 ;
      RECT 131.540000  62.135000 140.000000 112.450000 ;
    LAYER met4 ;
      RECT   0.000000   0.000000   1.670000   1.635000 ;
      RECT   0.000000   0.000000 140.000000   1.635000 ;
      RECT   0.000000   7.885000   1.670000   8.485000 ;
      RECT   0.000000   7.885000 140.000000   8.485000 ;
      RECT   0.000000  13.935000   1.365000  14.535000 ;
      RECT   0.000000  13.935000 140.000000  14.535000 ;
      RECT   0.000000  18.785000   1.365000  19.385000 ;
      RECT   0.000000  18.785000 140.000000  19.385000 ;
      RECT   0.000000  24.835000   1.670000  25.435000 ;
      RECT   0.000000  24.835000 140.000000  25.435000 ;
      RECT   0.000000  30.885000   1.670000  31.485000 ;
      RECT   0.000000  30.885000 140.000000  31.485000 ;
      RECT   0.000000  35.735000   1.670000  36.335000 ;
      RECT   0.000000  35.735000 140.000000  36.335000 ;
      RECT   0.000000  40.585000   1.670000  41.185000 ;
      RECT   0.000000  40.585000 140.000000  41.185000 ;
      RECT   0.000000  46.635000   1.670000  47.335000 ;
      RECT   0.000000  46.635000 140.000000  47.435000 ;
      RECT   0.000000  57.035000 140.000000  57.835000 ;
      RECT   0.000000  57.135000   1.670000  57.835000 ;
      RECT   0.000000  63.085000   1.670000  63.685000 ;
      RECT   0.000000  63.085000 140.000000  63.685000 ;
      RECT   0.000000  68.935000   1.670000  69.635000 ;
      RECT   0.000000  68.935000 140.000000  69.635000 ;
      RECT   0.000000  95.400000 140.000000 175.385000 ;
      RECT   1.365000  13.935000 138.635000  19.385000 ;
      RECT   1.365000  13.935000 138.635000  19.385000 ;
      RECT   1.570000  47.435000 138.430000  57.035000 ;
      RECT   1.670000   0.000000 137.855000 200.000000 ;
      RECT   1.670000   0.000000 138.330000   8.530000 ;
      RECT   1.670000   0.000000 138.330000   8.530000 ;
      RECT   1.670000   0.000000 138.330000   8.530000 ;
      RECT   1.670000   8.485000 140.000000   8.585000 ;
      RECT   1.670000   8.530000 137.855000  13.865000 ;
      RECT   1.670000   8.585000 138.430000   8.630000 ;
      RECT   1.670000   8.630000 137.955000  13.765000 ;
      RECT   1.670000  13.765000 138.430000  13.835000 ;
      RECT   1.670000  13.835000 140.000000  13.935000 ;
      RECT   1.670000  13.865000 138.330000  13.935000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  13.865000 138.330000 200.000000 ;
      RECT   1.670000  19.385000 138.330000  95.400000 ;
      RECT   1.670000 175.385000 138.330000 200.000000 ;
      RECT 138.330000   0.000000 140.000000   1.635000 ;
      RECT 138.330000   7.885000 140.000000   8.485000 ;
      RECT 138.330000  24.835000 140.000000  25.435000 ;
      RECT 138.330000  30.885000 140.000000  31.485000 ;
      RECT 138.330000  35.735000 140.000000  36.335000 ;
      RECT 138.330000  40.585000 140.000000  41.185000 ;
      RECT 138.330000  46.635000 140.000000  47.335000 ;
      RECT 138.330000  57.135000 140.000000  57.835000 ;
      RECT 138.330000  63.085000 140.000000  63.685000 ;
      RECT 138.330000  68.935000 140.000000  69.635000 ;
      RECT 138.635000  13.935000 140.000000  14.535000 ;
      RECT 138.635000  18.785000 140.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 140.000000   1.335000 ;
      RECT  0.000000  36.035000 140.000000  36.040000 ;
      RECT  0.000000  95.785000 140.000000 131.905000 ;
      RECT  0.000000 131.905000  39.295000 148.530000 ;
      RECT  0.000000 148.530000 140.000000 174.985000 ;
      RECT  1.765000  14.235000 138.235000  19.085000 ;
      RECT  2.070000   1.335000 137.930000  14.235000 ;
      RECT  2.070000  19.085000 137.930000  95.785000 ;
      RECT  2.070000 174.985000 137.930000 200.000000 ;
      RECT  9.605000  96.585000 126.350000 103.180000 ;
      RECT 11.565000 171.780000  99.610000 174.185000 ;
      RECT 63.935000 131.905000 140.000000 148.530000 ;
  END
END sky130_fd_io__top_gpio_ovtv2
END LIBRARY
