magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1217 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 493
rect 271 333 337 493
rect 439 333 505 493
rect 607 333 673 493
rect 879 333 945 493
rect 1047 333 1113 493
rect 103 289 1271 333
rect 22 215 340 255
rect 398 215 708 255
rect 770 215 1113 255
rect 1225 181 1271 289
rect 879 131 1271 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 18 289 69 527
rect 203 367 237 527
rect 371 367 405 527
rect 539 367 573 527
rect 707 367 845 527
rect 979 367 1013 527
rect 1147 367 1200 527
rect 18 147 757 181
rect 18 51 85 147
rect 119 17 153 113
rect 187 51 253 147
rect 355 131 421 147
rect 523 131 589 147
rect 691 131 757 147
rect 287 17 321 113
rect 439 51 1200 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 770 215 1113 255 6 A
port 1 nsew signal input
rlabel locali s 398 215 708 255 6 B
port 2 nsew signal input
rlabel locali s 22 215 340 255 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1217 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 879 131 1271 181 6 Y
port 8 nsew signal output
rlabel locali s 1225 181 1271 289 6 Y
port 8 nsew signal output
rlabel locali s 103 289 1271 333 6 Y
port 8 nsew signal output
rlabel locali s 1047 333 1113 493 6 Y
port 8 nsew signal output
rlabel locali s 879 333 945 493 6 Y
port 8 nsew signal output
rlabel locali s 607 333 673 493 6 Y
port 8 nsew signal output
rlabel locali s 439 333 505 493 6 Y
port 8 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 8 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1288 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1843154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1832018
<< end >>
