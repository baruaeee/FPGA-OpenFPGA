magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 544 157 827 203
rect 21 21 827 157
rect 29 -17 63 21
<< locali >>
rect 85 299 614 333
rect 657 299 723 493
rect 85 199 155 299
rect 483 283 614 299
rect 201 199 339 265
rect 373 199 431 265
rect 689 181 723 299
rect 657 51 723 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 401 123 493
rect 195 435 261 527
rect 351 401 417 493
rect 17 367 417 401
rect 507 367 572 527
rect 17 165 51 367
rect 757 299 811 527
rect 585 215 655 249
rect 585 165 621 215
rect 17 131 621 165
rect 17 56 105 131
rect 195 17 261 97
rect 351 51 417 131
rect 527 17 593 97
rect 757 17 811 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 201 199 339 265 6 A
port 1 nsew signal input
rlabel locali s 373 199 431 265 6 B
port 2 nsew signal input
rlabel locali s 483 283 614 299 6 C
port 3 nsew signal input
rlabel locali s 85 199 155 299 6 C
port 3 nsew signal input
rlabel locali s 85 299 614 333 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 21 21 827 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 544 157 827 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 657 51 723 181 6 X
port 8 nsew signal output
rlabel locali s 689 181 723 299 6 X
port 8 nsew signal output
rlabel locali s 657 299 723 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1660154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1653706
<< end >>
