magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 114 -17 148 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 835 47 865 177
rect 919 47 949 177
rect 1003 47 1033 177
rect 1087 47 1117 177
rect 1171 47 1201 177
rect 1255 47 1285 177
rect 1339 47 1369 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1003 297 1033 497
rect 1087 297 1117 497
rect 1171 297 1201 497
rect 1255 297 1285 497
rect 1339 297 1369 497
<< ndiff >>
rect 27 97 79 177
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 129 163 177
rect 109 95 119 129
rect 153 95 163 129
rect 109 47 163 95
rect 193 97 247 177
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 129 331 177
rect 277 95 287 129
rect 321 95 331 129
rect 277 47 331 95
rect 361 97 415 177
rect 361 63 371 97
rect 405 63 415 97
rect 361 47 415 63
rect 445 129 499 177
rect 445 95 455 129
rect 489 95 499 129
rect 445 47 499 95
rect 529 97 583 177
rect 529 63 539 97
rect 573 63 583 97
rect 529 47 583 63
rect 613 129 667 177
rect 613 95 623 129
rect 657 95 667 129
rect 613 47 667 95
rect 697 97 751 177
rect 697 63 707 97
rect 741 63 751 97
rect 697 47 751 63
rect 781 129 835 177
rect 781 95 791 129
rect 825 95 835 129
rect 781 47 835 95
rect 865 97 919 177
rect 865 63 875 97
rect 909 63 919 97
rect 865 47 919 63
rect 949 129 1003 177
rect 949 95 959 129
rect 993 95 1003 129
rect 949 47 1003 95
rect 1033 97 1087 177
rect 1033 63 1043 97
rect 1077 63 1087 97
rect 1033 47 1087 63
rect 1117 129 1171 177
rect 1117 95 1127 129
rect 1161 95 1171 129
rect 1117 47 1171 95
rect 1201 97 1255 177
rect 1201 63 1211 97
rect 1245 63 1255 97
rect 1201 47 1255 63
rect 1285 129 1339 177
rect 1285 95 1295 129
rect 1329 95 1339 129
rect 1285 47 1339 95
rect 1369 161 1445 177
rect 1369 127 1379 161
rect 1413 127 1445 161
rect 1369 93 1445 127
rect 1369 59 1379 93
rect 1413 59 1445 93
rect 1369 47 1445 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 479 163 497
rect 109 445 119 479
rect 153 445 163 479
rect 109 411 163 445
rect 109 377 119 411
rect 153 377 163 411
rect 109 343 163 377
rect 109 309 119 343
rect 153 309 163 343
rect 109 297 163 309
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 479 331 497
rect 277 445 287 479
rect 321 445 331 479
rect 277 411 331 445
rect 277 377 287 411
rect 321 377 331 411
rect 277 343 331 377
rect 277 309 287 343
rect 321 309 331 343
rect 277 297 331 309
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 463 499 497
rect 445 429 455 463
rect 489 429 499 463
rect 445 368 499 429
rect 445 334 455 368
rect 489 334 499 368
rect 445 297 499 334
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 463 667 497
rect 613 429 623 463
rect 657 429 667 463
rect 613 368 667 429
rect 613 334 623 368
rect 657 334 667 368
rect 613 297 667 334
rect 697 485 751 497
rect 697 451 707 485
rect 741 451 751 485
rect 697 417 751 451
rect 697 383 707 417
rect 741 383 751 417
rect 697 297 751 383
rect 781 463 835 497
rect 781 429 791 463
rect 825 429 835 463
rect 781 368 835 429
rect 781 334 791 368
rect 825 334 835 368
rect 781 297 835 334
rect 865 485 919 497
rect 865 451 875 485
rect 909 451 919 485
rect 865 417 919 451
rect 865 383 875 417
rect 909 383 919 417
rect 865 297 919 383
rect 949 463 1003 497
rect 949 429 959 463
rect 993 429 1003 463
rect 949 368 1003 429
rect 949 334 959 368
rect 993 334 1003 368
rect 949 297 1003 334
rect 1033 485 1087 497
rect 1033 451 1043 485
rect 1077 451 1087 485
rect 1033 417 1087 451
rect 1033 383 1043 417
rect 1077 383 1087 417
rect 1033 297 1087 383
rect 1117 463 1171 497
rect 1117 429 1127 463
rect 1161 429 1171 463
rect 1117 368 1171 429
rect 1117 334 1127 368
rect 1161 334 1171 368
rect 1117 297 1171 334
rect 1201 485 1255 497
rect 1201 451 1211 485
rect 1245 451 1255 485
rect 1201 417 1255 451
rect 1201 383 1211 417
rect 1245 383 1255 417
rect 1201 297 1255 383
rect 1285 463 1339 497
rect 1285 429 1295 463
rect 1329 429 1339 463
rect 1285 368 1339 429
rect 1285 334 1295 368
rect 1329 334 1339 368
rect 1285 297 1339 334
rect 1369 485 1445 497
rect 1369 451 1379 485
rect 1413 451 1445 485
rect 1369 417 1445 451
rect 1369 383 1379 417
rect 1413 383 1445 417
rect 1369 349 1445 383
rect 1369 315 1379 349
rect 1413 315 1445 349
rect 1369 297 1445 315
<< ndiffc >>
rect 35 63 69 97
rect 119 95 153 129
rect 203 63 237 97
rect 287 95 321 129
rect 371 63 405 97
rect 455 95 489 129
rect 539 63 573 97
rect 623 95 657 129
rect 707 63 741 97
rect 791 95 825 129
rect 875 63 909 97
rect 959 95 993 129
rect 1043 63 1077 97
rect 1127 95 1161 129
rect 1211 63 1245 97
rect 1295 95 1329 129
rect 1379 127 1413 161
rect 1379 59 1413 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 445 153 479
rect 119 377 153 411
rect 119 309 153 343
rect 203 451 237 485
rect 203 383 237 417
rect 287 445 321 479
rect 287 377 321 411
rect 287 309 321 343
rect 371 451 405 485
rect 371 383 405 417
rect 455 429 489 463
rect 455 334 489 368
rect 539 451 573 485
rect 539 383 573 417
rect 623 429 657 463
rect 623 334 657 368
rect 707 451 741 485
rect 707 383 741 417
rect 791 429 825 463
rect 791 334 825 368
rect 875 451 909 485
rect 875 383 909 417
rect 959 429 993 463
rect 959 334 993 368
rect 1043 451 1077 485
rect 1043 383 1077 417
rect 1127 429 1161 463
rect 1127 334 1161 368
rect 1211 451 1245 485
rect 1211 383 1245 417
rect 1295 429 1329 463
rect 1295 334 1329 368
rect 1379 451 1413 485
rect 1379 383 1413 417
rect 1379 315 1413 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1003 497 1033 523
rect 1087 497 1117 523
rect 1171 497 1201 523
rect 1255 497 1285 523
rect 1339 497 1369 523
rect 79 261 109 297
rect 27 259 109 261
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 27 249 361 259
rect 27 215 60 249
rect 94 215 128 249
rect 162 215 196 249
rect 230 215 264 249
rect 298 215 361 249
rect 27 205 361 215
rect 27 203 109 205
rect 79 177 109 203
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 751 259 781 297
rect 835 259 865 297
rect 919 259 949 297
rect 1003 259 1033 297
rect 1087 259 1117 297
rect 1171 259 1201 297
rect 1255 259 1285 297
rect 1339 259 1369 297
rect 415 249 1369 259
rect 415 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 707 249
rect 741 215 775 249
rect 809 215 843 249
rect 877 215 1369 249
rect 415 205 1369 215
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 751 177 781 205
rect 835 177 865 205
rect 919 177 949 205
rect 1003 177 1033 205
rect 1087 177 1117 205
rect 1171 177 1201 205
rect 1255 177 1285 205
rect 1339 177 1369 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 835 21 865 47
rect 919 21 949 47
rect 1003 21 1033 47
rect 1087 21 1117 47
rect 1171 21 1201 47
rect 1255 21 1285 47
rect 1339 21 1369 47
<< polycont >>
rect 60 215 94 249
rect 128 215 162 249
rect 196 215 230 249
rect 264 215 298 249
rect 435 215 469 249
rect 503 215 537 249
rect 571 215 605 249
rect 639 215 673 249
rect 707 215 741 249
rect 775 215 809 249
rect 843 215 877 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 367 69 383
rect 103 479 169 493
rect 103 445 119 479
rect 153 445 169 479
rect 103 411 169 445
rect 103 377 119 411
rect 153 377 169 411
rect 103 343 169 377
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 479 337 493
rect 271 445 287 479
rect 321 445 337 479
rect 271 411 337 445
rect 271 377 287 411
rect 321 377 337 411
rect 103 309 119 343
rect 153 323 169 343
rect 271 343 337 377
rect 371 485 405 527
rect 371 417 405 451
rect 371 367 405 383
rect 455 463 489 493
rect 455 368 489 429
rect 271 323 287 343
rect 153 309 287 323
rect 321 323 337 343
rect 523 485 589 527
rect 523 451 539 485
rect 573 451 589 485
rect 523 417 589 451
rect 523 383 539 417
rect 573 383 589 417
rect 523 367 589 383
rect 623 463 657 493
rect 623 368 657 429
rect 455 323 489 334
rect 691 485 757 527
rect 691 451 707 485
rect 741 451 757 485
rect 691 417 757 451
rect 691 383 707 417
rect 741 383 757 417
rect 691 367 757 383
rect 791 463 825 493
rect 791 368 825 429
rect 623 323 657 334
rect 859 485 925 527
rect 859 451 875 485
rect 909 451 925 485
rect 859 417 925 451
rect 859 383 875 417
rect 909 383 925 417
rect 859 367 925 383
rect 959 463 993 493
rect 959 368 993 429
rect 791 323 825 334
rect 1027 485 1093 527
rect 1027 451 1043 485
rect 1077 451 1093 485
rect 1027 417 1093 451
rect 1027 383 1043 417
rect 1077 383 1093 417
rect 1027 367 1093 383
rect 1127 463 1161 493
rect 1127 368 1161 429
rect 959 323 993 334
rect 1195 485 1261 527
rect 1195 451 1211 485
rect 1245 451 1261 485
rect 1195 417 1261 451
rect 1195 383 1211 417
rect 1245 383 1261 417
rect 1195 367 1261 383
rect 1295 463 1329 493
rect 1295 368 1329 429
rect 1127 323 1161 334
rect 1295 323 1329 334
rect 321 309 403 323
rect 103 289 403 309
rect 455 289 1329 323
rect 1363 485 1429 527
rect 1363 451 1379 485
rect 1413 451 1429 485
rect 1363 417 1429 451
rect 1363 383 1379 417
rect 1413 383 1429 417
rect 1363 349 1429 383
rect 1363 315 1379 349
rect 1413 315 1429 349
rect 1363 297 1429 315
rect 27 249 332 255
rect 27 215 60 249
rect 94 215 128 249
rect 162 215 196 249
rect 230 215 264 249
rect 298 215 332 249
rect 368 249 403 289
rect 368 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 707 249
rect 741 215 775 249
rect 809 215 843 249
rect 877 215 893 249
rect 368 181 403 215
rect 942 181 1329 289
rect 119 147 403 181
rect 455 147 1329 181
rect 119 129 153 147
rect 19 97 85 113
rect 19 63 35 97
rect 69 63 85 97
rect 19 17 85 63
rect 287 129 321 147
rect 119 51 153 95
rect 187 97 253 113
rect 187 63 203 97
rect 237 63 253 97
rect 187 17 253 63
rect 455 129 489 147
rect 287 52 321 95
rect 355 97 421 113
rect 355 63 371 97
rect 405 63 421 97
rect 355 17 421 63
rect 623 129 657 147
rect 455 51 489 95
rect 523 97 589 113
rect 523 63 539 97
rect 573 63 589 97
rect 523 17 589 63
rect 791 129 825 147
rect 623 51 657 95
rect 691 97 757 113
rect 691 63 707 97
rect 741 63 757 97
rect 691 17 757 63
rect 959 129 993 147
rect 791 51 825 95
rect 859 97 925 113
rect 859 63 875 97
rect 909 63 925 97
rect 859 17 925 63
rect 1127 129 1161 147
rect 959 51 993 95
rect 1027 97 1093 113
rect 1027 63 1043 97
rect 1077 63 1093 97
rect 1027 17 1093 63
rect 1295 129 1329 147
rect 1127 51 1161 95
rect 1195 97 1261 113
rect 1195 63 1211 97
rect 1245 63 1261 97
rect 1195 17 1261 63
rect 1295 51 1329 95
rect 1363 161 1429 177
rect 1363 127 1379 161
rect 1413 127 1429 161
rect 1363 93 1429 127
rect 1363 59 1379 93
rect 1413 59 1429 93
rect 1363 17 1429 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 298 221 332 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 942 153 976 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 942 221 976 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 206 221 240 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 114 -17 148 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 114 527 148 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 942 289 976 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 114 221 148 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 46 221 80 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 114 527 148 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 114 -17 148 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 114 -17 148 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 114 527 148 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 buf_12
rlabel metal1 s 0 -48 1472 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 3147130
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3135996
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
