magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 35 21 643 203
rect 35 17 64 21
rect 30 -17 64 17
<< locali >>
rect 111 165 157 493
rect 293 199 358 282
rect 111 127 191 165
rect 153 51 191 127
rect 448 73 524 265
rect 562 150 625 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 333 77 527
rect 191 444 257 527
rect 295 384 358 493
rect 191 338 358 384
rect 392 387 437 493
rect 471 425 537 527
rect 571 387 615 493
rect 191 199 259 338
rect 392 334 615 387
rect 225 165 259 199
rect 225 131 373 165
rect 53 17 119 93
rect 225 17 291 89
rect 335 51 373 131
rect 561 17 627 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 448 73 524 265 6 A1
port 1 nsew signal input
rlabel locali s 562 150 625 265 6 A2
port 2 nsew signal input
rlabel locali s 293 199 358 282 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 35 17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 35 21 643 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 153 51 191 127 6 X
port 8 nsew signal output
rlabel locali s 111 127 191 165 6 X
port 8 nsew signal output
rlabel locali s 111 165 157 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4102614
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4097060
<< end >>
