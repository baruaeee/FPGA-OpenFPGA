magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 21 1839 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 776 47 806 177
rect 860 47 890 177
rect 1053 47 1083 177
rect 1137 47 1167 177
rect 1211 47 1241 177
rect 1295 47 1325 177
rect 1379 47 1409 177
rect 1479 47 1509 177
rect 1563 47 1593 177
rect 1647 47 1677 177
rect 1731 47 1761 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 514 297 544 497
rect 598 297 628 497
rect 687 297 717 497
rect 776 297 806 497
rect 860 297 890 497
rect 1005 297 1035 497
rect 1127 297 1157 497
rect 1211 297 1241 497
rect 1295 297 1325 497
rect 1379 297 1409 497
rect 1479 297 1509 497
rect 1563 297 1593 497
rect 1647 297 1677 497
rect 1731 297 1761 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 97 163 131
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 161 247 177
rect 193 127 203 161
rect 237 127 247 161
rect 193 93 247 127
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 97 331 131
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 161 413 177
rect 361 127 371 161
rect 405 127 413 161
rect 361 93 413 127
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 467 95 519 177
rect 467 61 475 95
rect 509 61 519 95
rect 467 47 519 61
rect 549 163 603 177
rect 549 129 559 163
rect 593 129 603 163
rect 549 47 603 129
rect 633 119 687 177
rect 633 85 643 119
rect 677 85 687 119
rect 633 47 687 85
rect 717 93 776 177
rect 717 59 729 93
rect 763 59 776 93
rect 717 47 776 59
rect 806 119 860 177
rect 806 85 816 119
rect 850 85 860 119
rect 806 47 860 85
rect 890 93 942 177
rect 890 59 900 93
rect 934 59 942 93
rect 890 47 942 59
rect 996 101 1053 177
rect 996 67 1004 101
rect 1038 67 1053 101
rect 996 47 1053 67
rect 1083 93 1137 177
rect 1083 59 1093 93
rect 1127 59 1137 93
rect 1083 47 1137 59
rect 1167 47 1211 177
rect 1241 93 1295 177
rect 1241 59 1251 93
rect 1285 59 1295 93
rect 1241 47 1295 59
rect 1325 47 1379 177
rect 1409 93 1479 177
rect 1409 59 1427 93
rect 1461 59 1479 93
rect 1409 47 1479 59
rect 1509 131 1563 177
rect 1509 97 1519 131
rect 1553 97 1563 131
rect 1509 47 1563 97
rect 1593 97 1647 177
rect 1593 63 1603 97
rect 1637 63 1647 97
rect 1593 47 1647 63
rect 1677 131 1731 177
rect 1677 97 1687 131
rect 1721 97 1731 131
rect 1677 47 1731 97
rect 1761 161 1813 177
rect 1761 127 1771 161
rect 1805 127 1813 161
rect 1761 93 1813 127
rect 1761 59 1771 93
rect 1805 59 1813 93
rect 1761 47 1813 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 483 163 497
rect 109 449 119 483
rect 153 449 163 483
rect 109 415 163 449
rect 109 381 119 415
rect 153 381 163 415
rect 109 347 163 381
rect 109 313 119 347
rect 153 313 163 347
rect 109 297 163 313
rect 193 489 247 497
rect 193 455 203 489
rect 237 455 247 489
rect 193 421 247 455
rect 193 387 203 421
rect 237 387 247 421
rect 193 353 247 387
rect 193 319 203 353
rect 237 319 247 353
rect 193 297 247 319
rect 277 483 331 497
rect 277 449 287 483
rect 321 449 331 483
rect 277 415 331 449
rect 277 381 287 415
rect 321 381 331 415
rect 277 347 331 381
rect 277 313 287 347
rect 321 313 331 347
rect 277 297 331 313
rect 361 485 514 497
rect 361 315 371 485
rect 473 315 514 485
rect 361 297 514 315
rect 544 455 598 497
rect 544 421 554 455
rect 588 421 598 455
rect 544 387 598 421
rect 544 353 554 387
rect 588 353 598 387
rect 544 297 598 353
rect 628 471 687 497
rect 628 437 638 471
rect 672 437 687 471
rect 628 297 687 437
rect 717 297 776 497
rect 806 475 860 497
rect 806 441 816 475
rect 850 441 860 475
rect 806 297 860 441
rect 890 297 1005 497
rect 1035 475 1127 497
rect 1035 441 1064 475
rect 1098 441 1127 475
rect 1035 297 1127 441
rect 1157 455 1211 497
rect 1157 421 1167 455
rect 1201 421 1211 455
rect 1157 297 1211 421
rect 1241 475 1295 497
rect 1241 441 1251 475
rect 1285 441 1295 475
rect 1241 297 1295 441
rect 1325 455 1379 497
rect 1325 421 1335 455
rect 1369 421 1379 455
rect 1325 297 1379 421
rect 1409 475 1479 497
rect 1409 441 1427 475
rect 1461 441 1479 475
rect 1409 297 1479 441
rect 1509 467 1563 497
rect 1509 433 1519 467
rect 1553 433 1563 467
rect 1509 359 1563 433
rect 1509 325 1519 359
rect 1553 325 1563 359
rect 1509 297 1563 325
rect 1593 485 1647 497
rect 1593 451 1603 485
rect 1637 451 1647 485
rect 1593 401 1647 451
rect 1593 367 1603 401
rect 1637 367 1647 401
rect 1593 297 1647 367
rect 1677 467 1731 497
rect 1677 433 1687 467
rect 1721 433 1731 467
rect 1677 359 1731 433
rect 1677 325 1687 359
rect 1721 325 1731 359
rect 1677 297 1731 325
rect 1761 485 1813 497
rect 1761 451 1771 485
rect 1805 451 1813 485
rect 1761 417 1813 451
rect 1761 383 1771 417
rect 1805 383 1813 417
rect 1761 349 1813 383
rect 1761 315 1771 349
rect 1805 315 1813 349
rect 1761 297 1813 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 131 153 165
rect 119 63 153 97
rect 203 127 237 161
rect 203 59 237 93
rect 287 131 321 165
rect 287 63 321 97
rect 371 127 405 161
rect 371 59 405 93
rect 475 61 509 95
rect 559 129 593 163
rect 643 85 677 119
rect 729 59 763 93
rect 816 85 850 119
rect 900 59 934 93
rect 1004 67 1038 101
rect 1093 59 1127 93
rect 1251 59 1285 93
rect 1427 59 1461 93
rect 1519 97 1553 131
rect 1603 63 1637 97
rect 1687 97 1721 131
rect 1771 127 1805 161
rect 1771 59 1805 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 449 153 483
rect 119 381 153 415
rect 119 313 153 347
rect 203 455 237 489
rect 203 387 237 421
rect 203 319 237 353
rect 287 449 321 483
rect 287 381 321 415
rect 287 313 321 347
rect 371 315 473 485
rect 554 421 588 455
rect 554 353 588 387
rect 638 437 672 471
rect 816 441 850 475
rect 1064 441 1098 475
rect 1167 421 1201 455
rect 1251 441 1285 475
rect 1335 421 1369 455
rect 1427 441 1461 475
rect 1519 433 1553 467
rect 1519 325 1553 359
rect 1603 451 1637 485
rect 1603 367 1637 401
rect 1687 433 1721 467
rect 1687 325 1721 359
rect 1771 451 1805 485
rect 1771 383 1805 417
rect 1771 315 1805 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 514 497 544 523
rect 598 497 628 523
rect 687 497 717 523
rect 776 497 806 523
rect 860 497 890 523
rect 1005 497 1035 523
rect 1127 497 1157 523
rect 1211 497 1241 523
rect 1295 497 1325 523
rect 1379 497 1409 523
rect 1479 497 1509 523
rect 1563 497 1593 523
rect 1647 497 1677 523
rect 1731 497 1761 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 514 265 544 297
rect 598 265 628 297
rect 687 265 717 297
rect 776 265 806 297
rect 860 265 890 297
rect 1005 265 1035 297
rect 1127 265 1157 297
rect 1211 265 1241 297
rect 1295 265 1325 297
rect 1379 265 1409 297
rect 1479 265 1509 297
rect 1563 265 1593 297
rect 1647 265 1677 297
rect 1731 265 1761 297
rect 79 249 472 265
rect 79 215 360 249
rect 394 215 428 249
rect 462 215 472 249
rect 79 199 472 215
rect 514 249 633 265
rect 514 215 584 249
rect 618 215 633 249
rect 514 199 633 215
rect 675 249 729 265
rect 675 215 685 249
rect 719 215 729 249
rect 675 199 729 215
rect 776 249 963 265
rect 776 215 910 249
rect 944 215 963 249
rect 1005 249 1169 265
rect 1005 235 1125 249
rect 776 199 963 215
rect 1043 215 1125 235
rect 1159 215 1169 249
rect 1043 199 1169 215
rect 1211 249 1325 265
rect 1211 215 1229 249
rect 1263 215 1325 249
rect 1211 199 1325 215
rect 1367 249 1421 265
rect 1367 215 1377 249
rect 1411 215 1421 249
rect 1367 199 1421 215
rect 1479 249 1761 265
rect 1479 215 1527 249
rect 1561 215 1595 249
rect 1629 215 1761 249
rect 1479 199 1761 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 519 177 549 199
rect 603 177 633 199
rect 687 177 717 199
rect 776 177 806 199
rect 860 177 890 199
rect 1053 177 1083 199
rect 1137 177 1167 199
rect 1211 177 1241 199
rect 1295 177 1325 199
rect 1379 177 1409 199
rect 1479 177 1509 199
rect 1563 177 1593 199
rect 1647 177 1677 199
rect 1731 177 1761 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 776 21 806 47
rect 860 21 890 47
rect 1053 21 1083 47
rect 1137 21 1167 47
rect 1211 21 1241 47
rect 1295 21 1325 47
rect 1379 21 1409 47
rect 1479 21 1509 47
rect 1563 21 1593 47
rect 1647 21 1677 47
rect 1731 21 1761 47
<< polycont >>
rect 360 215 394 249
rect 428 215 462 249
rect 584 215 618 249
rect 685 215 719 249
rect 910 215 944 249
rect 1125 215 1159 249
rect 1229 215 1263 249
rect 1377 215 1411 249
rect 1527 215 1561 249
rect 1595 215 1629 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 27 485 69 527
rect 27 451 35 485
rect 203 489 237 527
rect 27 417 69 451
rect 27 383 35 417
rect 27 349 69 383
rect 27 315 35 349
rect 27 299 69 315
rect 103 449 119 483
rect 153 449 169 483
rect 103 415 169 449
rect 103 381 119 415
rect 153 381 169 415
rect 103 347 169 381
rect 103 313 119 347
rect 153 313 169 347
rect 103 267 169 313
rect 371 485 473 527
rect 203 421 237 455
rect 203 353 237 387
rect 203 303 237 319
rect 271 449 287 483
rect 321 449 337 483
rect 271 415 337 449
rect 271 381 287 415
rect 321 381 337 415
rect 271 347 337 381
rect 271 313 287 347
rect 321 313 337 347
rect 638 471 672 527
rect 1048 475 1114 527
rect 554 455 588 471
rect 638 421 672 437
rect 706 441 816 475
rect 850 441 866 475
rect 1048 441 1064 475
rect 1098 441 1114 475
rect 1235 475 1301 527
rect 1167 455 1201 471
rect 554 387 588 421
rect 706 387 740 441
rect 1235 441 1251 475
rect 1285 441 1301 475
rect 1411 475 1477 527
rect 1587 485 1645 527
rect 1335 455 1369 471
rect 1167 405 1201 421
rect 1411 441 1427 475
rect 1461 441 1477 475
rect 1519 467 1553 483
rect 1335 405 1369 421
rect 271 267 310 313
rect 371 299 473 315
rect 516 353 554 387
rect 588 353 740 387
rect 774 371 1479 405
rect 103 213 310 267
rect 516 249 550 353
rect 774 319 808 371
rect 344 215 360 249
rect 394 215 428 249
rect 462 215 550 249
rect 27 161 69 177
rect 27 127 35 161
rect 27 93 69 127
rect 27 59 35 93
rect 103 165 169 213
rect 103 131 119 165
rect 153 131 169 165
rect 103 97 169 131
rect 103 63 119 97
rect 153 63 169 97
rect 203 161 237 177
rect 203 93 237 127
rect 27 17 69 59
rect 271 165 310 213
rect 271 131 287 165
rect 321 131 337 165
rect 271 97 337 131
rect 271 63 287 97
rect 321 63 337 97
rect 371 161 419 177
rect 405 127 419 161
rect 516 163 550 215
rect 584 285 808 319
rect 842 301 1362 335
rect 584 249 618 285
rect 842 249 876 301
rect 664 215 685 249
rect 719 215 876 249
rect 910 249 944 265
rect 1125 249 1159 301
rect 1316 265 1362 301
rect 944 215 1091 233
rect 584 199 618 215
rect 910 199 1091 215
rect 1125 199 1159 215
rect 1217 249 1263 265
rect 1217 215 1229 249
rect 1057 175 1091 199
rect 1057 169 1099 175
rect 1057 165 1107 169
rect 1217 165 1263 215
rect 1316 249 1411 265
rect 1316 215 1377 249
rect 1316 199 1411 215
rect 1445 249 1479 371
rect 1519 359 1553 433
rect 1587 451 1603 485
rect 1637 451 1645 485
rect 1771 485 1813 527
rect 1587 401 1645 451
rect 1587 367 1603 401
rect 1637 367 1645 401
rect 1587 351 1645 367
rect 1681 467 1737 483
rect 1681 433 1687 467
rect 1721 433 1737 467
rect 1681 359 1737 433
rect 1519 317 1553 325
rect 1681 325 1687 359
rect 1721 325 1737 359
rect 1681 317 1737 325
rect 1519 283 1737 317
rect 1805 451 1813 485
rect 1771 417 1813 451
rect 1805 383 1813 417
rect 1771 349 1813 383
rect 1805 315 1813 349
rect 1771 299 1813 315
rect 1445 215 1527 249
rect 1561 215 1595 249
rect 1629 215 1645 249
rect 516 129 559 163
rect 593 129 609 163
rect 643 129 1023 163
rect 1057 146 1263 165
rect 1445 163 1479 215
rect 1681 181 1737 283
rect 1059 144 1263 146
rect 1062 142 1263 144
rect 1064 139 1263 142
rect 1067 135 1263 139
rect 1069 131 1263 135
rect 371 93 419 127
rect 643 119 677 129
rect 203 17 237 59
rect 405 59 419 93
rect 454 61 475 95
rect 509 85 643 95
rect 816 119 850 129
rect 509 61 677 85
rect 371 17 419 59
rect 711 59 729 93
rect 763 59 782 93
rect 984 117 1023 129
rect 1341 129 1479 163
rect 1519 147 1737 181
rect 1519 131 1569 147
rect 984 101 1038 117
rect 816 69 850 85
rect 711 17 782 59
rect 884 59 900 93
rect 934 59 950 93
rect 884 17 950 59
rect 984 67 1004 101
rect 1341 93 1375 129
rect 1553 97 1569 131
rect 1681 131 1737 147
rect 984 51 1038 67
rect 1077 59 1093 93
rect 1127 59 1143 93
rect 1235 59 1251 93
rect 1285 59 1375 93
rect 1411 59 1427 93
rect 1461 59 1477 93
rect 1519 63 1569 97
rect 1603 97 1645 113
rect 1637 63 1645 97
rect 1681 97 1687 131
rect 1721 97 1737 131
rect 1681 63 1737 97
rect 1771 161 1813 177
rect 1805 127 1813 161
rect 1771 93 1813 127
rect 1077 17 1143 59
rect 1411 17 1477 59
rect 1603 17 1645 63
rect 1805 59 1813 93
rect 1771 17 1813 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 1316 221 1350 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1684 357 1718 391 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 1684 85 1718 119 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 122 85 156 119 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 122 357 156 391 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 122 425 156 459 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 1684 425 1718 459 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 1316 289 1350 323 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1224 221 1258 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1224 153 1258 187 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1684 153 1718 187 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 1684 221 1718 255 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 1684 289 1718 323 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
rlabel comment s 0 0 0 0 4 ha_4
rlabel metal1 s 0 -48 1840 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1840 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_END 2190846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2176828
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 46.000 0.000 
<< end >>
