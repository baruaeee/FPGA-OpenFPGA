/home/exotic/Desktop/FPGA-OpenFPGA/PNR/auto_3x3_sky_scl/lef/IO/sky130_fd_io__corner_bus_overlay.lef