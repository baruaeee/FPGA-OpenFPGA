VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
  MACRO oaTaper STRING ;
END PROPERTYDEFINITIONS

MACRO DFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX1 0 0 ;
  SIZE 9.2 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.787937 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 0.385 1.05 1.625 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 8.585 2.44 8.87 3.45 ;
        RECT 8.61 0.68 8.87 3.45 ;
        RECT 8.585 0.68 8.87 1.33 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 7.69 2.44 7.955 3.45 ;
        RECT 7.69 0.68 7.955 1.33 ;
        RECT 7.69 0.68 7.95 3.45 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER met1 ;
      ANTENNAMAXAREACAR 2.620159 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 2.974603 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 6.77 1.405 7.03 2.645 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.91746 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.079365 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 2.315 1.05 3.555 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 9.2 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 9.2 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 6.345 0.765 6.575 3.53 ;
      RECT 5.915 0.765 6.575 0.995 ;
      RECT 5.915 0.705 6.145 0.995 ;
      RECT 1.435 3.375 3.905 3.605 ;
      RECT 3.675 2.505 3.905 3.605 ;
      RECT 1.435 0.705 1.665 3.605 ;
      RECT 2.725 2.945 2.955 3.235 ;
      RECT 1.865 2.945 2.095 3.235 ;
      RECT 1.865 3.005 2.955 3.175 ;
      RECT 7.205 0.61 7.435 3.53 ;
      RECT 4.965 1.145 5.195 2.795 ;
      RECT 4.535 0.705 4.765 3.235 ;
      RECT 4.105 0.705 4.335 3.235 ;
      RECT 3.245 0.705 3.475 3.235 ;
      RECT 0.145 0.705 0.375 3.235 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END DFFRX1

MACRO TBUFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1 0 0 ;
  SIZE 3.68 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 3.09 2.52 3.535 3.53 ;
        RECT 3.09 0.61 3.535 1.26 ;
        RECT 3.09 0.61 3.35 3.53 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 3.68 0.2 ;
    END
  END VSS
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER met1 ;
      ANTENNAMAXAREACAR 1.370794 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.504762 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 1.85 1.05 3.09 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER met1 ;
      ANTENNAMAXAREACAR 0.86619 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.911111 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.71 1.665 1.97 2.905 ;
    END
  END A
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 3.68 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 2.385 3.24 2.615 3.53 ;
      RECT 2.43 0.785 2.57 3.53 ;
      RECT 2.385 1.82 2.615 2.11 ;
      RECT 2.375 0.785 2.605 1.075 ;
      RECT 1.435 3.24 1.665 3.53 ;
      RECT 1.43 0.685 1.57 3.385 ;
      RECT 1.34 1.48 1.57 1.77 ;
      RECT 1.005 0.61 1.235 0.9 ;
      RECT 1.005 0.685 1.62 0.825 ;
      RECT 0.145 3.24 0.375 3.53 ;
      RECT 0.175 0.61 0.345 3.53 ;
      RECT 0.145 1.82 0.375 2.11 ;
      RECT 0.145 0.61 0.375 0.9 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END TBUFX1

MACRO CLKINVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX1 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.545 2.905 1.05 3.495 ;
        RECT 0.79 0.64 1.05 3.495 ;
        RECT 0.545 0.64 1.05 0.87 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2835 LAYER met1 ;
      ANTENNAMAXAREACAR 0.308818 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.33 1.19 0.59 2.43 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END CLKINVX1

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.575 2.84 1.05 3.49 ;
        RECT 0.79 0.605 1.05 3.49 ;
        RECT 0.575 0.605 1.05 1.255 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2835 LAYER met1 ;
      ANTENNAMAXAREACAR 0.308818 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.33 1.43 0.59 2.67 ;
    END
  END A
END INVX1

MACRO MX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X1 0 0 ;
  SIZE 3.68 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 2.755 2.91 3.35 3.5 ;
        RECT 3.09 0.64 3.35 3.5 ;
        RECT 2.755 0.64 3.35 1.23 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.555873 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.653968 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 0.48 1.05 1.72 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER met1 ;
      ANTENNAMAXAREACAR 2.112857 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 2.060317 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 2.28 1.05 3.52 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.674603 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.793651 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 2.17 0.875 2.43 2.115 ;
    END
  END B
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 3.68 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 3.68 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 1.435 0.655 1.665 3.38 ;
      RECT 1.435 2.29 2.84 2.52 ;
      RECT 2.61 2 2.84 2.52 ;
      RECT 0.145 0.655 0.375 3.38 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END MX2X1

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 2.3 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.78254 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.920635 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 1.455 1.05 2.695 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 2.3 0.2 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.593651 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.698413 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.33 1.145 0.59 2.385 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.495 3.21 1.97 3.5 ;
        RECT 1.71 0.505 1.97 3.5 ;
        RECT 1.495 0.505 1.97 0.795 ;
    END
  END Y
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 2.3 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 0.115 3.27 1.2 3.5 ;
      RECT 0.97 2.84 1.2 3.5 ;
      RECT 1.19 0.965 1.42 3.07 ;
      RECT 0.765 0.965 1.42 1.195 ;
      RECT 0.765 0.475 0.995 1.195 ;
      RECT 0.545 0.475 0.995 0.705 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END OR2X1

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 2.3 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 2.3 0.2 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5292 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.065 3.23 1.51 3.52 ;
        RECT 1.25 0.61 1.51 3.52 ;
        RECT 1.065 0.61 1.51 1.26 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.949841 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.11746 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 1.685 1.05 2.925 ;
    END
  END A
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 2.3 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 0.145 3.24 0.375 3.53 ;
      RECT 0.145 0.655 0.285 3.53 ;
      RECT 0.145 1.48 0.515 1.77 ;
      RECT 0.145 0.655 0.375 0.945 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END BUFX2

MACRO CLKAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X2 0 0 ;
  SIZE 2.3 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 2.3 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 2.3 4.34 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5292 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.49 3.24 1.97 3.53 ;
        RECT 1.71 0.68 1.97 3.53 ;
        RECT 1.495 0.68 1.97 1.33 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22125 LAYER met1 ;
      ANTENNAMAXAREACAR 0.718418 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.845198 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.25 1.685 1.51 2.925 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22125 LAYER met1 ;
      ANTENNAMAXAREACAR 0.537853 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.632768 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.33 1.855 0.59 3.095 ;
    END
  END B
  OBS
    LAYER met1 ;
      RECT 0.575 3.24 0.96 3.53 ;
      RECT 0.73 1.55 0.96 3.53 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END CLKAND2X2

MACRO DFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX1 0 0 ;
  SIZE 11.5 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 10.245 2.42 10.71 3.57 ;
        RECT 10.45 0.57 10.71 3.57 ;
        RECT 10.245 0.57 10.71 1.35 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.50085 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 10.91 2.42 11.275 3.57 ;
        RECT 10.91 0.57 11.275 1.35 ;
        RECT 10.91 0.57 11.17 3.57 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 11.5 0.2 ;
    END
  END VSS
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER met1 ;
      ANTENNAMAXAREACAR 1.75127 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.952381 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 4.01 1.075 4.27 2.315 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 1.009206 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.187302 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 2.19 1.05 3.43 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.868889 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.022222 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 6.77 1.155 7.03 2.395 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.631429 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.742857 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 0.805 1.05 2.045 ;
    END
  END D
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 11.5 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 5.945 0.845 8.545 1.015 ;
      RECT 8.315 0.705 8.545 1.015 ;
      RECT 5.945 0.705 6.175 1.015 ;
      RECT 5.555 3.425 8.545 3.595 ;
      RECT 8.315 3.26 8.545 3.595 ;
      RECT 5.555 3.26 5.785 3.595 ;
      RECT 5.125 2.535 5.355 3.235 ;
      RECT 5.125 2.535 8.38 2.765 ;
      RECT 5.515 0.705 5.745 2.765 ;
      RECT 7.885 2.945 8.115 3.235 ;
      RECT 6.415 2.945 6.645 3.235 ;
      RECT 6.415 3.005 8.115 3.175 ;
      RECT 3.405 3.005 4.925 3.235 ;
      RECT 4.695 0.715 4.925 3.235 ;
      RECT 3.405 2.945 3.635 3.235 ;
      RECT 4.695 0.715 5.315 0.945 ;
      RECT 5.085 0.655 5.315 0.945 ;
      RECT 1.435 3.405 3.265 3.575 ;
      RECT 3.095 2.165 3.265 3.575 ;
      RECT 1.435 0.705 1.665 3.575 ;
      RECT 3.095 2.165 3.325 2.455 ;
      RECT 9.695 0.705 9.925 3.235 ;
      RECT 8.835 0.705 9.065 3.235 ;
      RECT 6.345 0.535 8.145 0.705 ;
      RECT 3.215 0.715 4.365 0.885 ;
      RECT 2.725 0.705 2.955 3.235 ;
      RECT 0.145 0.705 0.375 3.235 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END DFFSRX1

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 1.84 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5178 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.575 3.21 1.51 3.47 ;
        RECT 1.25 0.655 1.51 3.47 ;
        RECT 0.975 0.655 1.51 0.915 ;
        RECT 0.575 2.82 0.805 3.47 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2835 LAYER met1 ;
      ANTENNAMAXAREACAR 0.428748 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.504409 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.33 1.29 0.59 2.53 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2835 LAYER met1 ;
      ANTENNAMAXAREACAR 0.437743 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.514991 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 1.19 1.05 2.43 ;
    END
  END B
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.84 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.84 4.34 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END NAND2X1

MACRO CLKBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX2 0 0 ;
  SIZE 2.3 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 2.3 0.2 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5292 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.065 3.24 1.51 3.53 ;
        RECT 1.25 0.61 1.51 3.53 ;
        RECT 1.065 0.61 1.51 1.26 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.949841 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.11746 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 1.805 1.05 3.045 ;
    END
  END A
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 2.3 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 0.145 3.24 0.375 3.53 ;
      RECT 0.145 0.655 0.285 3.53 ;
      RECT 0.145 1.48 0.375 1.77 ;
      RECT 0.145 0.655 0.375 0.945 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END CLKBUFX2

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.567 LAYER met1 ;
      ANTENNAMAXAREACAR 0.376279 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.382716 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.33 1.29 0.59 2.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5292 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.575 2.735 1.05 3.385 ;
        RECT 0.79 0.61 1.05 3.385 ;
        RECT 0.575 0.61 1.05 0.9 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
    END
  END VDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END INVX2

MACRO CLKMX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X2 0 0 ;
  SIZE 3.68 BY 4.14 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.315 LAYER met1 ;
      ANTENNAMAXAREACAR 1.08746 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 1.095238 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 1.25 1.69 1.51 2.93 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.787937 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 0.79 2.02 1.05 3.26 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER met1 ;
      ANTENNAMAXAREACAR 0.771746 LAYER met1 ;
      ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 2.17 1.505 2.43 2.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5292 LAYER met1 ;
    PORT
      LAYER met1 ;
        RECT 2.63 0.68 3.015 3.45 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 3.68 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 3.68 4.34 ;
    END
  END VDD
  OBS
    LAYER met1 ;
      RECT 1.435 3.24 1.88 3.53 ;
      RECT 1.65 0.705 1.88 3.53 ;
      RECT 1.435 0.705 1.88 0.995 ;
      RECT 0.145 0.705 0.375 3.235 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END CLKMX2X2

END LIBRARY
