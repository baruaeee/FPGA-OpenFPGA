magic
tech sky130A
magscale 1 2
timestamp 1729530005
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 183
rect 29 -17 63 21
<< scnmos >>
rect 79 47 657 157
<< scpmoshvt >>
rect 79 323 657 497
<< ndiff >>
rect 27 112 79 157
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 657 112 709 157
rect 657 78 667 112
rect 701 78 709 112
rect 657 47 709 78
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 383 79 451
rect 27 349 35 383
rect 69 349 79 383
rect 27 323 79 349
rect 657 485 709 497
rect 657 451 667 485
rect 701 451 709 485
rect 657 383 709 451
rect 657 349 667 383
rect 701 349 709 383
rect 657 323 709 349
<< ndiffc >>
rect 35 78 69 112
rect 667 78 701 112
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 667 451 701 485
rect 667 349 701 383
<< poly >>
rect 79 497 657 523
rect 79 297 657 323
rect 79 275 343 297
rect 79 241 95 275
rect 129 241 194 275
rect 228 241 293 275
rect 327 241 343 275
rect 79 225 343 241
rect 385 239 657 255
rect 385 205 401 239
rect 435 205 504 239
rect 538 205 607 239
rect 641 205 657 239
rect 385 183 657 205
rect 79 157 657 183
rect 79 21 657 47
<< polycont >>
rect 95 241 129 275
rect 194 241 228 275
rect 293 241 327 275
rect 401 205 435 239
rect 504 205 538 239
rect 607 205 641 239
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 485 719 493
rect 17 459 35 485
rect 69 459 667 485
rect 701 459 719 485
rect 17 425 29 459
rect 69 451 121 459
rect 63 425 121 451
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 397 459
rect 431 425 489 459
rect 523 425 581 459
rect 615 451 667 459
rect 615 425 673 451
rect 707 425 719 459
rect 17 383 719 425
rect 17 349 35 383
rect 69 349 667 383
rect 701 349 719 383
rect 17 309 719 349
rect 17 241 95 275
rect 129 241 194 275
rect 228 241 293 275
rect 327 241 347 275
rect 17 171 347 241
rect 381 239 719 309
rect 381 205 401 239
rect 435 205 504 239
rect 538 205 607 239
rect 641 205 719 239
rect 17 112 719 171
rect 17 78 35 112
rect 69 78 667 112
rect 701 78 719 112
rect 17 17 719 78
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 451 35 459
rect 35 451 63 459
rect 29 425 63 451
rect 121 425 155 459
rect 213 425 247 459
rect 305 425 339 459
rect 397 425 431 459
rect 489 425 523 459
rect 581 425 615 459
rect 673 451 701 459
rect 701 451 707 459
rect 673 425 707 451
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 14 459 722 468
rect 14 428 29 459
rect 17 425 29 428
rect 63 425 121 459
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 397 459
rect 431 425 489 459
rect 523 425 581 459
rect 615 425 673 459
rect 707 428 722 459
rect 707 425 719 428
rect 17 416 719 425
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 33 429 68 460 0 FreeSans 200 0 0 0 KAPWR
port 1 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 lpflow_decapkapwr_8
rlabel metal1 s 17 416 719 428 1 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 722 468 1 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -48 736 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 2334036
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2329784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
