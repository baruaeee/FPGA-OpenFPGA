/home/exotic/Desktop/FPGA-OpenFPGA/PNR/auto_3x3_gpdk/lef/gsclib045_lvt_macro.lef