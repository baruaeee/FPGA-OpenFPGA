/home/exotic/Desktop/FPGA-OpenFPGA/PNR/auto_3x3_sky_scl/lef/IO/sky130_fd_io__top_power_hvc_wpadv2.lef